// *!***************************************************************************
// *! Copyright 2019 International Business Machines
// *!
// *! Licensed under the Apache License, Version 2.0 (the "License");
// *! you may not use this file except in compliance with the License.
// *! You may obtain a copy of the License at
// *! http://www.apache.org/licenses/LICENSE-2.0
// *!
// *! The patent license granted to you in Section 3 of the License, as applied
// *! to the "Work," hereby includes implementations of the Work in physical form.
// *!
// *! Unless required by applicable law or agreed to in writing, the reference design
// *! distributed under the License is distributed on an "AS IS" BASIS,
// *! WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// *! See the License for the specific language governing permissions and
// *! limitations under the License.
// *!
// *! The background Specification upon which this is based is managed by and available from
// *! the OpenCAPI Consortium.  More information can be found at https://opencapi.org.
// *!***************************************************************************
 
`timescale 1ns / 1ps

 


module ocx_dlx_crc (

    init                     // < input 
  , checkbits_in             // < input 
  , data                     // < input 
  , checkbits0_out            // > output  
  , checkbits1_out

);

input           init;
input  [35:0]   checkbits_in;
input  [511:0]  data;
output [35:0]   checkbits0_out;
output [35:0]   checkbits1_out;

wire [35:0]  checkbits,temp_checkbits0, temp_checkbits1;
//wire [0:511] dat;



assign  checkbits = init ? 36'b0 : checkbits_in;



assign temp_checkbits0[35] = checkbits[1] ^ checkbits[3] ^ checkbits[4] ^ checkbits[5] ^ checkbits[7] ^ checkbits[8] ^ checkbits[10] ^ checkbits[11] ^ checkbits[12] ^ checkbits[14] ^ checkbits[15] ^ checkbits[17] ^ checkbits[19] ^ checkbits[22] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[29] ^ checkbits[30] ^ checkbits[31] ^ checkbits[32] ^ data[2] ^ data[3] ^ data[5] ^ data[8] ^ data[10] ^ data[12] ^ data[13] ^ data[15] ^ data[17] ^ data[18] ^ data[19] ^ data[21] ^ data[22] ^ data[23] ^ data[25] ^ data[31] ^ data[33] ^ data[35] ^ data[37] ^ data[38] ^ data[41] ^ data[43] ^ data[46] ^ data[49] ^ data[50] ^ data[52] ^ data[55] ^ data[57] ^ data[59] ^ data[61] ^ data[62] ^ data[63] ^ data[64] ^ data[66] ^ data[68] ^ data[69] ^ data[77] ^ data[81] ^ data[85] ^ data[86] ^ data[93] ^ data[95] ^ data[97] ^ data[98] ^ data[99] ^ data[100] ^ data[102] ^ data[103] ^ data[104] ^ data[105] ^ data[107] ^ data[108] ^ data[111] ^ data[112] ^ data[119] ^ data[120] ^ data[122] ^ data[123] ^ data[124] ^ data[127] ^ data[130] ^ data[132] ^ data[134] ^ data[135] ^ data[136] ^ data[137] ^ data[138] ^ data[139] ^ data[141] ^ data[142] ^ data[143] ^ data[146] ^ data[148] ^ data[151] ^ data[153] ^ data[154] ^ data[155] ^ data[156] ^ data[157] ^ data[158] ^ data[166] ^ data[167] ^ data[168] ^ data[170] ^ data[171] ^ data[172] ^ data[176] ^ data[177] ^ data[178] ^ data[182] ^ data[183] ^ data[188] ^ data[192] ^ data[194] ^ data[195] ^ data[196] ^ data[197] ^ data[199] ^ data[204] ^ data[207] ^ data[210] ^ data[211] ^ data[218] ^ data[219] ^ data[220] ^ data[222] ^ data[223] ^ data[225] ^ data[226] ^ data[232] ^ data[233] ^ data[235] ^ data[239] ^ data[241] ^ data[242] ^ data[244] ^ data[245] ^ data[246] ^ data[247] ^ data[251] ^ data[252] ^ data[253] ;

assign temp_checkbits0[34] = checkbits[0] ^ checkbits[2] ^ checkbits[3] ^ checkbits[4] ^ checkbits[6] ^ checkbits[7] ^ checkbits[9] ^ checkbits[10] ^ checkbits[11] ^ checkbits[13] ^ checkbits[14] ^ checkbits[16] ^ checkbits[18] ^ checkbits[21] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[29] ^ checkbits[30] ^ checkbits[31] ^ data[3] ^ data[4] ^ data[6] ^ data[9] ^ data[11] ^ data[13] ^ data[14] ^ data[16] ^ data[18] ^ data[19] ^ data[20] ^ data[22] ^ data[23] ^ data[24] ^ data[26] ^ data[32] ^ data[34] ^ data[36] ^ data[38] ^ data[39] ^ data[42] ^ data[44] ^ data[47] ^ data[50] ^ data[51] ^ data[53] ^ data[56] ^ data[58] ^ data[60] ^ data[62] ^ data[63] ^ data[64] ^ data[65] ^ data[67] ^ data[69] ^ data[70] ^ data[78] ^ data[82] ^ data[86] ^ data[87] ^ data[94] ^ data[96] ^ data[98] ^ data[99] ^ data[100] ^ data[101] ^ data[103] ^ data[104] ^ data[105] ^ data[106] ^ data[108] ^ data[109] ^ data[112] ^ data[113] ^ data[120] ^ data[121] ^ data[123] ^ data[124] ^ data[125] ^ data[128] ^ data[131] ^ data[133] ^ data[135] ^ data[136] ^ data[137] ^ data[138] ^ data[139] ^ data[140] ^ data[142] ^ data[143] ^ data[144] ^ data[147] ^ data[149] ^ data[152] ^ data[154] ^ data[155] ^ data[156] ^ data[157] ^ data[158] ^ data[159] ^ data[167] ^ data[168] ^ data[169] ^ data[171] ^ data[172] ^ data[173] ^ data[177] ^ data[178] ^ data[179] ^ data[183] ^ data[184] ^ data[189] ^ data[193] ^ data[195] ^ data[196] ^ data[197] ^ data[198] ^ data[200] ^ data[205] ^ data[208] ^ data[211] ^ data[212] ^ data[219] ^ data[220] ^ data[221] ^ data[223] ^ data[224] ^ data[226] ^ data[227] ^ data[233] ^ data[234] ^ data[236] ^ data[240] ^ data[242] ^ data[243] ^ data[245] ^ data[246] ^ data[247] ^ data[248] ^ data[252] ^ data[253] ^ data[254] ;

assign temp_checkbits0[33] = checkbits[2] ^ checkbits[4] ^ checkbits[6] ^ checkbits[7] ^ checkbits[9] ^ checkbits[11] ^ checkbits[13] ^ checkbits[14] ^ checkbits[19] ^ checkbits[20] ^ checkbits[22] ^ checkbits[23] ^ checkbits[24] ^ checkbits[31] ^ checkbits[32] ^ data[0] ^ data[2] ^ data[3] ^ data[4] ^ data[7] ^ data[8] ^ data[13] ^ data[14] ^ data[18] ^ data[20] ^ data[22] ^ data[24] ^ data[27] ^ data[31] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[45] ^ data[46] ^ data[48] ^ data[49] ^ data[50] ^ data[51] ^ data[54] ^ data[55] ^ data[62] ^ data[65] ^ data[69] ^ data[70] ^ data[71] ^ data[77] ^ data[79] ^ data[81] ^ data[83] ^ data[85] ^ data[86] ^ data[87] ^ data[88] ^ data[93] ^ data[98] ^ data[101] ^ data[103] ^ data[106] ^ data[108] ^ data[109] ^ data[110] ^ data[111] ^ data[112] ^ data[113] ^ data[114] ^ data[119] ^ data[120] ^ data[121] ^ data[123] ^ data[125] ^ data[126] ^ data[127] ^ data[129] ^ data[130] ^ data[135] ^ data[140] ^ data[142] ^ data[144] ^ data[145] ^ data[146] ^ data[150] ^ data[151] ^ data[154] ^ data[159] ^ data[160] ^ data[166] ^ data[167] ^ data[169] ^ data[171] ^ data[173] ^ data[174] ^ data[176] ^ data[177] ^ data[179] ^ data[180] ^ data[182] ^ data[183] ^ data[184] ^ data[185] ^ data[188] ^ data[190] ^ data[192] ^ data[195] ^ data[198] ^ data[201] ^ data[204] ^ data[206] ^ data[207] ^ data[209] ^ data[210] ^ data[211] ^ data[212] ^ data[213] ^ data[218] ^ data[219] ^ data[221] ^ data[223] ^ data[224] ^ data[226] ^ data[227] ^ data[228] ^ data[232] ^ data[233] ^ data[234] ^ data[237] ^ data[239] ^ data[242] ^ data[243] ^ data[245] ^ data[248] ^ data[249] ^ data[251] ^ data[252] ^ data[254] ^ data[255] ;

assign temp_checkbits0[32] = checkbits[1] ^ checkbits[3] ^ checkbits[5] ^ checkbits[6] ^ checkbits[8] ^ checkbits[10] ^ checkbits[12] ^ checkbits[13] ^ checkbits[18] ^ checkbits[19] ^ checkbits[21] ^ checkbits[22] ^ checkbits[23] ^ checkbits[30] ^ checkbits[31] ^ checkbits[35] ^ data[1] ^ data[3] ^ data[4] ^ data[5] ^ data[8] ^ data[9] ^ data[14] ^ data[15] ^ data[19] ^ data[21] ^ data[23] ^ data[25] ^ data[28] ^ data[32] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[46] ^ data[47] ^ data[49] ^ data[50] ^ data[51] ^ data[52] ^ data[55] ^ data[56] ^ data[63] ^ data[66] ^ data[70] ^ data[71] ^ data[72] ^ data[78] ^ data[80] ^ data[82] ^ data[84] ^ data[86] ^ data[87] ^ data[88] ^ data[89] ^ data[94] ^ data[99] ^ data[102] ^ data[104] ^ data[107] ^ data[109] ^ data[110] ^ data[111] ^ data[112] ^ data[113] ^ data[114] ^ data[115] ^ data[120] ^ data[121] ^ data[122] ^ data[124] ^ data[126] ^ data[127] ^ data[128] ^ data[130] ^ data[131] ^ data[136] ^ data[141] ^ data[143] ^ data[145] ^ data[146] ^ data[147] ^ data[151] ^ data[152] ^ data[155] ^ data[160] ^ data[161] ^ data[167] ^ data[168] ^ data[170] ^ data[172] ^ data[174] ^ data[175] ^ data[177] ^ data[178] ^ data[180] ^ data[181] ^ data[183] ^ data[184] ^ data[185] ^ data[186] ^ data[189] ^ data[191] ^ data[193] ^ data[196] ^ data[199] ^ data[202] ^ data[205] ^ data[207] ^ data[208] ^ data[210] ^ data[211] ^ data[212] ^ data[213] ^ data[214] ^ data[219] ^ data[220] ^ data[222] ^ data[224] ^ data[225] ^ data[227] ^ data[228] ^ data[229] ^ data[233] ^ data[234] ^ data[235] ^ data[238] ^ data[240] ^ data[243] ^ data[244] ^ data[246] ^ data[249] ^ data[250] ^ data[252] ^ data[253] ^ data[255] ;

assign temp_checkbits0[31] = checkbits[0] ^ checkbits[2] ^ checkbits[4] ^ checkbits[5] ^ checkbits[7] ^ checkbits[9] ^ checkbits[11] ^ checkbits[12] ^ checkbits[17] ^ checkbits[18] ^ checkbits[20] ^ checkbits[21] ^ checkbits[22] ^ checkbits[29] ^ checkbits[30] ^ checkbits[34] ^ checkbits[35] ^ data[2] ^ data[4] ^ data[5] ^ data[6] ^ data[9] ^ data[10] ^ data[15] ^ data[16] ^ data[20] ^ data[22] ^ data[24] ^ data[26] ^ data[29] ^ data[33] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[47] ^ data[48] ^ data[50] ^ data[51] ^ data[52] ^ data[53] ^ data[56] ^ data[57] ^ data[64] ^ data[67] ^ data[71] ^ data[72] ^ data[73] ^ data[79] ^ data[81] ^ data[83] ^ data[85] ^ data[87] ^ data[88] ^ data[89] ^ data[90] ^ data[95] ^ data[100] ^ data[103] ^ data[105] ^ data[108] ^ data[110] ^ data[111] ^ data[112] ^ data[113] ^ data[114] ^ data[115] ^ data[116] ^ data[121] ^ data[122] ^ data[123] ^ data[125] ^ data[127] ^ data[128] ^ data[129] ^ data[131] ^ data[132] ^ data[137] ^ data[142] ^ data[144] ^ data[146] ^ data[147] ^ data[148] ^ data[152] ^ data[153] ^ data[156] ^ data[161] ^ data[162] ^ data[168] ^ data[169] ^ data[171] ^ data[173] ^ data[175] ^ data[176] ^ data[178] ^ data[179] ^ data[181] ^ data[182] ^ data[184] ^ data[185] ^ data[186] ^ data[187] ^ data[190] ^ data[192] ^ data[194] ^ data[197] ^ data[200] ^ data[203] ^ data[206] ^ data[208] ^ data[209] ^ data[211] ^ data[212] ^ data[213] ^ data[214] ^ data[215] ^ data[220] ^ data[221] ^ data[223] ^ data[225] ^ data[226] ^ data[228] ^ data[229] ^ data[230] ^ data[234] ^ data[235] ^ data[236] ^ data[239] ^ data[241] ^ data[244] ^ data[245] ^ data[247] ^ data[250] ^ data[251] ^ data[253] ^ data[254] ;

assign temp_checkbits0[30] = checkbits[5] ^ checkbits[6] ^ checkbits[7] ^ checkbits[12] ^ checkbits[14] ^ checkbits[15] ^ checkbits[16] ^ checkbits[20] ^ checkbits[21] ^ checkbits[22] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[30] ^ checkbits[31] ^ checkbits[32] ^ checkbits[33] ^ checkbits[34] ^ data[0] ^ data[2] ^ data[6] ^ data[7] ^ data[8] ^ data[11] ^ data[12] ^ data[13] ^ data[15] ^ data[16] ^ data[18] ^ data[19] ^ data[22] ^ data[27] ^ data[30] ^ data[31] ^ data[33] ^ data[34] ^ data[35] ^ data[37] ^ data[38] ^ data[42] ^ data[44] ^ data[46] ^ data[48] ^ data[50] ^ data[51] ^ data[53] ^ data[54] ^ data[55] ^ data[58] ^ data[59] ^ data[61] ^ data[62] ^ data[63] ^ data[64] ^ data[65] ^ data[66] ^ data[69] ^ data[72] ^ data[73] ^ data[74] ^ data[77] ^ data[80] ^ data[81] ^ data[82] ^ data[84] ^ data[85] ^ data[88] ^ data[89] ^ data[90] ^ data[91] ^ data[93] ^ data[95] ^ data[96] ^ data[97] ^ data[98] ^ data[99] ^ data[100] ^ data[101] ^ data[102] ^ data[103] ^ data[105] ^ data[106] ^ data[107] ^ data[108] ^ data[109] ^ data[113] ^ data[114] ^ data[115] ^ data[116] ^ data[117] ^ data[119] ^ data[120] ^ data[126] ^ data[127] ^ data[128] ^ data[129] ^ data[133] ^ data[134] ^ data[135] ^ data[136] ^ data[137] ^ data[139] ^ data[141] ^ data[142] ^ data[145] ^ data[146] ^ data[147] ^ data[149] ^ data[151] ^ data[155] ^ data[156] ^ data[158] ^ data[162] ^ data[163] ^ data[166] ^ data[167] ^ data[168] ^ data[169] ^ data[171] ^ data[174] ^ data[178] ^ data[179] ^ data[180] ^ data[185] ^ data[186] ^ data[187] ^ data[191] ^ data[192] ^ data[193] ^ data[194] ^ data[196] ^ data[197] ^ data[198] ^ data[199] ^ data[201] ^ data[209] ^ data[211] ^ data[212] ^ data[213] ^ data[214] ^ data[215] ^ data[216] ^ data[218] ^ data[219] ^ data[220] ^ data[221] ^ data[223] ^ data[224] ^ data[225] ^ data[227] ^ data[229] ^ data[230] ^ data[231] ^ data[232] ^ data[233] ^ data[236] ^ data[237] ^ data[239] ^ data[240] ^ data[241] ^ data[244] ^ data[247] ^ data[248] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[29] = checkbits[1] ^ checkbits[3] ^ checkbits[6] ^ checkbits[7] ^ checkbits[8] ^ checkbits[10] ^ checkbits[12] ^ checkbits[13] ^ checkbits[17] ^ checkbits[20] ^ checkbits[21] ^ checkbits[22] ^ checkbits[24] ^ checkbits[27] ^ checkbits[28] ^ checkbits[33] ^ data[1] ^ data[2] ^ data[5] ^ data[7] ^ data[9] ^ data[10] ^ data[14] ^ data[15] ^ data[16] ^ data[18] ^ data[20] ^ data[21] ^ data[22] ^ data[25] ^ data[28] ^ data[32] ^ data[33] ^ data[34] ^ data[36] ^ data[37] ^ data[39] ^ data[41] ^ data[45] ^ data[46] ^ data[47] ^ data[50] ^ data[51] ^ data[54] ^ data[56] ^ data[57] ^ data[60] ^ data[61] ^ data[65] ^ data[67] ^ data[68] ^ data[69] ^ data[70] ^ data[73] ^ data[74] ^ data[75] ^ data[77] ^ data[78] ^ data[82] ^ data[83] ^ data[89] ^ data[90] ^ data[91] ^ data[92] ^ data[93] ^ data[94] ^ data[95] ^ data[96] ^ data[101] ^ data[105] ^ data[106] ^ data[109] ^ data[110] ^ data[111] ^ data[112] ^ data[114] ^ data[115] ^ data[116] ^ data[117] ^ data[118] ^ data[119] ^ data[121] ^ data[122] ^ data[123] ^ data[124] ^ data[128] ^ data[129] ^ data[132] ^ data[139] ^ data[140] ^ data[141] ^ data[147] ^ data[150] ^ data[151] ^ data[152] ^ data[153] ^ data[154] ^ data[155] ^ data[158] ^ data[159] ^ data[163] ^ data[164] ^ data[166] ^ data[169] ^ data[171] ^ data[175] ^ data[176] ^ data[177] ^ data[178] ^ data[179] ^ data[180] ^ data[181] ^ data[182] ^ data[183] ^ data[186] ^ data[187] ^ data[193] ^ data[196] ^ data[198] ^ data[200] ^ data[202] ^ data[204] ^ data[207] ^ data[211] ^ data[212] ^ data[213] ^ data[214] ^ data[215] ^ data[216] ^ data[217] ^ data[218] ^ data[221] ^ data[223] ^ data[224] ^ data[228] ^ data[230] ^ data[231] ^ data[234] ^ data[235] ^ data[237] ^ data[238] ^ data[239] ^ data[240] ^ data[244] ^ data[246] ^ data[247] ^ data[248] ^ data[249] ^ data[251] ^ data[252] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[28] = checkbits[0] ^ checkbits[2] ^ checkbits[5] ^ checkbits[6] ^ checkbits[7] ^ checkbits[9] ^ checkbits[11] ^ checkbits[12] ^ checkbits[16] ^ checkbits[19] ^ checkbits[20] ^ checkbits[21] ^ checkbits[23] ^ checkbits[26] ^ checkbits[27] ^ checkbits[32] ^ checkbits[35] ^ data[2] ^ data[3] ^ data[6] ^ data[8] ^ data[10] ^ data[11] ^ data[15] ^ data[16] ^ data[17] ^ data[19] ^ data[21] ^ data[22] ^ data[23] ^ data[26] ^ data[29] ^ data[33] ^ data[34] ^ data[35] ^ data[37] ^ data[38] ^ data[40] ^ data[42] ^ data[46] ^ data[47] ^ data[48] ^ data[51] ^ data[52] ^ data[55] ^ data[57] ^ data[58] ^ data[61] ^ data[62] ^ data[66] ^ data[68] ^ data[69] ^ data[70] ^ data[71] ^ data[74] ^ data[75] ^ data[76] ^ data[78] ^ data[79] ^ data[83] ^ data[84] ^ data[90] ^ data[91] ^ data[92] ^ data[93] ^ data[94] ^ data[95] ^ data[96] ^ data[97] ^ data[102] ^ data[106] ^ data[107] ^ data[110] ^ data[111] ^ data[112] ^ data[113] ^ data[115] ^ data[116] ^ data[117] ^ data[118] ^ data[119] ^ data[120] ^ data[122] ^ data[123] ^ data[124] ^ data[125] ^ data[129] ^ data[130] ^ data[133] ^ data[140] ^ data[141] ^ data[142] ^ data[148] ^ data[151] ^ data[152] ^ data[153] ^ data[154] ^ data[155] ^ data[156] ^ data[159] ^ data[160] ^ data[164] ^ data[165] ^ data[167] ^ data[170] ^ data[172] ^ data[176] ^ data[177] ^ data[178] ^ data[179] ^ data[180] ^ data[181] ^ data[182] ^ data[183] ^ data[184] ^ data[187] ^ data[188] ^ data[194] ^ data[197] ^ data[199] ^ data[201] ^ data[203] ^ data[205] ^ data[208] ^ data[212] ^ data[213] ^ data[214] ^ data[215] ^ data[216] ^ data[217] ^ data[218] ^ data[219] ^ data[222] ^ data[224] ^ data[225] ^ data[229] ^ data[231] ^ data[232] ^ data[235] ^ data[236] ^ data[238] ^ data[239] ^ data[240] ^ data[241] ^ data[245] ^ data[247] ^ data[248] ^ data[249] ^ data[250] ^ data[252] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[27] = checkbits[1] ^ checkbits[4] ^ checkbits[5] ^ checkbits[6] ^ checkbits[8] ^ checkbits[10] ^ checkbits[11] ^ checkbits[15] ^ checkbits[18] ^ checkbits[19] ^ checkbits[20] ^ checkbits[22] ^ checkbits[25] ^ checkbits[26] ^ checkbits[31] ^ checkbits[34] ^ data[0] ^ data[3] ^ data[4] ^ data[7] ^ data[9] ^ data[11] ^ data[12] ^ data[16] ^ data[17] ^ data[18] ^ data[20] ^ data[22] ^ data[23] ^ data[24] ^ data[27] ^ data[30] ^ data[34] ^ data[35] ^ data[36] ^ data[38] ^ data[39] ^ data[41] ^ data[43] ^ data[47] ^ data[48] ^ data[49] ^ data[52] ^ data[53] ^ data[56] ^ data[58] ^ data[59] ^ data[62] ^ data[63] ^ data[67] ^ data[69] ^ data[70] ^ data[71] ^ data[72] ^ data[75] ^ data[76] ^ data[77] ^ data[79] ^ data[80] ^ data[84] ^ data[85] ^ data[91] ^ data[92] ^ data[93] ^ data[94] ^ data[95] ^ data[96] ^ data[97] ^ data[98] ^ data[103] ^ data[107] ^ data[108] ^ data[111] ^ data[112] ^ data[113] ^ data[114] ^ data[116] ^ data[117] ^ data[118] ^ data[119] ^ data[120] ^ data[121] ^ data[123] ^ data[124] ^ data[125] ^ data[126] ^ data[130] ^ data[131] ^ data[134] ^ data[141] ^ data[142] ^ data[143] ^ data[149] ^ data[152] ^ data[153] ^ data[154] ^ data[155] ^ data[156] ^ data[157] ^ data[160] ^ data[161] ^ data[165] ^ data[166] ^ data[168] ^ data[171] ^ data[173] ^ data[177] ^ data[178] ^ data[179] ^ data[180] ^ data[181] ^ data[182] ^ data[183] ^ data[184] ^ data[185] ^ data[188] ^ data[189] ^ data[195] ^ data[198] ^ data[200] ^ data[202] ^ data[204] ^ data[206] ^ data[209] ^ data[213] ^ data[214] ^ data[215] ^ data[216] ^ data[217] ^ data[218] ^ data[219] ^ data[220] ^ data[223] ^ data[225] ^ data[226] ^ data[230] ^ data[232] ^ data[233] ^ data[236] ^ data[237] ^ data[239] ^ data[240] ^ data[241] ^ data[242] ^ data[246] ^ data[248] ^ data[249] ^ data[250] ^ data[251] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[26] = checkbits[0] ^ checkbits[1] ^ checkbits[8] ^ checkbits[9] ^ checkbits[11] ^ checkbits[12] ^ checkbits[15] ^ checkbits[18] ^ checkbits[21] ^ checkbits[22] ^ checkbits[24] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[29] ^ checkbits[31] ^ checkbits[32] ^ checkbits[33] ^ checkbits[35] ^ data[1] ^ data[2] ^ data[3] ^ data[4] ^ data[15] ^ data[22] ^ data[24] ^ data[28] ^ data[33] ^ data[36] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[46] ^ data[48] ^ data[52] ^ data[53] ^ data[54] ^ data[55] ^ data[60] ^ data[61] ^ data[62] ^ data[66] ^ data[69] ^ data[70] ^ data[71] ^ data[72] ^ data[73] ^ data[76] ^ data[78] ^ data[80] ^ data[92] ^ data[94] ^ data[96] ^ data[100] ^ data[102] ^ data[103] ^ data[105] ^ data[107] ^ data[109] ^ data[111] ^ data[113] ^ data[114] ^ data[115] ^ data[117] ^ data[118] ^ data[121] ^ data[123] ^ data[125] ^ data[126] ^ data[130] ^ data[131] ^ data[134] ^ data[136] ^ data[137] ^ data[138] ^ data[139] ^ data[141] ^ data[144] ^ data[146] ^ data[148] ^ data[150] ^ data[151] ^ data[161] ^ data[162] ^ data[168] ^ data[169] ^ data[170] ^ data[171] ^ data[174] ^ data[176] ^ data[177] ^ data[179] ^ data[180] ^ data[181] ^ data[184] ^ data[185] ^ data[186] ^ data[188] ^ data[189] ^ data[190] ^ data[192] ^ data[194] ^ data[195] ^ data[197] ^ data[201] ^ data[203] ^ data[204] ^ data[205] ^ data[211] ^ data[214] ^ data[215] ^ data[216] ^ data[217] ^ data[221] ^ data[222] ^ data[223] ^ data[224] ^ data[225] ^ data[227] ^ data[231] ^ data[232] ^ data[234] ^ data[235] ^ data[237] ^ data[238] ^ data[239] ^ data[240] ^ data[243] ^ data[244] ^ data[245] ^ data[246] ^ data[249] ^ data[250] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[25] = checkbits[0] ^ checkbits[7] ^ checkbits[8] ^ checkbits[10] ^ checkbits[11] ^ checkbits[14] ^ checkbits[17] ^ checkbits[20] ^ checkbits[21] ^ checkbits[23] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[30] ^ checkbits[31] ^ checkbits[32] ^ checkbits[34] ^ data[0] ^ data[2] ^ data[3] ^ data[4] ^ data[5] ^ data[16] ^ data[23] ^ data[25] ^ data[29] ^ data[34] ^ data[37] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[47] ^ data[49] ^ data[53] ^ data[54] ^ data[55] ^ data[56] ^ data[61] ^ data[62] ^ data[63] ^ data[67] ^ data[70] ^ data[71] ^ data[72] ^ data[73] ^ data[74] ^ data[77] ^ data[79] ^ data[81] ^ data[93] ^ data[95] ^ data[97] ^ data[101] ^ data[103] ^ data[104] ^ data[106] ^ data[108] ^ data[110] ^ data[112] ^ data[114] ^ data[115] ^ data[116] ^ data[118] ^ data[119] ^ data[122] ^ data[124] ^ data[126] ^ data[127] ^ data[131] ^ data[132] ^ data[135] ^ data[137] ^ data[138] ^ data[139] ^ data[140] ^ data[142] ^ data[145] ^ data[147] ^ data[149] ^ data[151] ^ data[152] ^ data[162] ^ data[163] ^ data[169] ^ data[170] ^ data[171] ^ data[172] ^ data[175] ^ data[177] ^ data[178] ^ data[180] ^ data[181] ^ data[182] ^ data[185] ^ data[186] ^ data[187] ^ data[189] ^ data[190] ^ data[191] ^ data[193] ^ data[195] ^ data[196] ^ data[198] ^ data[202] ^ data[204] ^ data[205] ^ data[206] ^ data[212] ^ data[215] ^ data[216] ^ data[217] ^ data[218] ^ data[222] ^ data[223] ^ data[224] ^ data[225] ^ data[226] ^ data[228] ^ data[232] ^ data[233] ^ data[235] ^ data[236] ^ data[238] ^ data[239] ^ data[240] ^ data[241] ^ data[244] ^ data[245] ^ data[246] ^ data[247] ^ data[250] ^ data[251] ^ data[254] ^ data[255] ;

assign temp_checkbits0[24] = checkbits[6] ^ checkbits[7] ^ checkbits[9] ^ checkbits[10] ^ checkbits[13] ^ checkbits[16] ^ checkbits[19] ^ checkbits[20] ^ checkbits[22] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[29] ^ checkbits[30] ^ checkbits[31] ^ checkbits[33] ^ checkbits[35] ^ data[0] ^ data[1] ^ data[3] ^ data[4] ^ data[5] ^ data[6] ^ data[17] ^ data[24] ^ data[26] ^ data[30] ^ data[35] ^ data[38] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[46] ^ data[48] ^ data[50] ^ data[54] ^ data[55] ^ data[56] ^ data[57] ^ data[62] ^ data[63] ^ data[64] ^ data[68] ^ data[71] ^ data[72] ^ data[73] ^ data[74] ^ data[75] ^ data[78] ^ data[80] ^ data[82] ^ data[94] ^ data[96] ^ data[98] ^ data[102] ^ data[104] ^ data[105] ^ data[107] ^ data[109] ^ data[111] ^ data[113] ^ data[115] ^ data[116] ^ data[117] ^ data[119] ^ data[120] ^ data[123] ^ data[125] ^ data[127] ^ data[128] ^ data[132] ^ data[133] ^ data[136] ^ data[138] ^ data[139] ^ data[140] ^ data[141] ^ data[143] ^ data[146] ^ data[148] ^ data[150] ^ data[152] ^ data[153] ^ data[163] ^ data[164] ^ data[170] ^ data[171] ^ data[172] ^ data[173] ^ data[176] ^ data[178] ^ data[179] ^ data[181] ^ data[182] ^ data[183] ^ data[186] ^ data[187] ^ data[188] ^ data[190] ^ data[191] ^ data[192] ^ data[194] ^ data[196] ^ data[197] ^ data[199] ^ data[203] ^ data[205] ^ data[206] ^ data[207] ^ data[213] ^ data[216] ^ data[217] ^ data[218] ^ data[219] ^ data[223] ^ data[224] ^ data[225] ^ data[226] ^ data[227] ^ data[229] ^ data[233] ^ data[234] ^ data[236] ^ data[237] ^ data[239] ^ data[240] ^ data[241] ^ data[242] ^ data[245] ^ data[246] ^ data[247] ^ data[248] ^ data[251] ^ data[252] ^ data[255] ;

assign temp_checkbits0[23] = checkbits[1] ^ checkbits[3] ^ checkbits[4] ^ checkbits[6] ^ checkbits[7] ^ checkbits[9] ^ checkbits[10] ^ checkbits[11] ^ checkbits[14] ^ checkbits[17] ^ checkbits[18] ^ checkbits[21] ^ checkbits[22] ^ checkbits[23] ^ checkbits[24] ^ checkbits[27] ^ checkbits[31] ^ checkbits[34] ^ checkbits[35] ^ data[1] ^ data[3] ^ data[4] ^ data[6] ^ data[7] ^ data[8] ^ data[10] ^ data[12] ^ data[13] ^ data[15] ^ data[17] ^ data[19] ^ data[21] ^ data[22] ^ data[23] ^ data[27] ^ data[33] ^ data[35] ^ data[36] ^ data[37] ^ data[38] ^ data[39] ^ data[42] ^ data[44] ^ data[45] ^ data[47] ^ data[50] ^ data[51] ^ data[52] ^ data[56] ^ data[58] ^ data[59] ^ data[61] ^ data[62] ^ data[65] ^ data[66] ^ data[68] ^ data[72] ^ data[73] ^ data[74] ^ data[75] ^ data[76] ^ data[77] ^ data[79] ^ data[83] ^ data[85] ^ data[86] ^ data[93] ^ data[98] ^ data[100] ^ data[102] ^ data[104] ^ data[106] ^ data[107] ^ data[110] ^ data[111] ^ data[114] ^ data[116] ^ data[117] ^ data[118] ^ data[119] ^ data[121] ^ data[122] ^ data[123] ^ data[126] ^ data[127] ^ data[128] ^ data[129] ^ data[130] ^ data[132] ^ data[133] ^ data[135] ^ data[136] ^ data[138] ^ data[140] ^ data[143] ^ data[144] ^ data[146] ^ data[147] ^ data[148] ^ data[149] ^ data[155] ^ data[156] ^ data[157] ^ data[158] ^ data[164] ^ data[165] ^ data[166] ^ data[167] ^ data[168] ^ data[170] ^ data[173] ^ data[174] ^ data[176] ^ data[178] ^ data[179] ^ data[180] ^ data[184] ^ data[187] ^ data[189] ^ data[191] ^ data[193] ^ data[194] ^ data[196] ^ data[198] ^ data[199] ^ data[200] ^ data[206] ^ data[208] ^ data[210] ^ data[211] ^ data[214] ^ data[217] ^ data[222] ^ data[223] ^ data[224] ^ data[227] ^ data[228] ^ data[230] ^ data[232] ^ data[233] ^ data[234] ^ data[237] ^ data[238] ^ data[239] ^ data[240] ^ data[243] ^ data[244] ^ data[245] ^ data[248] ^ data[249] ^ data[251] ;

assign temp_checkbits0[22] = checkbits[0] ^ checkbits[2] ^ checkbits[3] ^ checkbits[5] ^ checkbits[6] ^ checkbits[8] ^ checkbits[9] ^ checkbits[10] ^ checkbits[13] ^ checkbits[16] ^ checkbits[17] ^ checkbits[20] ^ checkbits[21] ^ checkbits[22] ^ checkbits[23] ^ checkbits[26] ^ checkbits[30] ^ checkbits[33] ^ checkbits[34] ^ data[2] ^ data[4] ^ data[5] ^ data[7] ^ data[8] ^ data[9] ^ data[11] ^ data[13] ^ data[14] ^ data[16] ^ data[18] ^ data[20] ^ data[22] ^ data[23] ^ data[24] ^ data[28] ^ data[34] ^ data[36] ^ data[37] ^ data[38] ^ data[39] ^ data[40] ^ data[43] ^ data[45] ^ data[46] ^ data[48] ^ data[51] ^ data[52] ^ data[53] ^ data[57] ^ data[59] ^ data[60] ^ data[62] ^ data[63] ^ data[66] ^ data[67] ^ data[69] ^ data[73] ^ data[74] ^ data[75] ^ data[76] ^ data[77] ^ data[78] ^ data[80] ^ data[84] ^ data[86] ^ data[87] ^ data[94] ^ data[99] ^ data[101] ^ data[103] ^ data[105] ^ data[107] ^ data[108] ^ data[111] ^ data[112] ^ data[115] ^ data[117] ^ data[118] ^ data[119] ^ data[120] ^ data[122] ^ data[123] ^ data[124] ^ data[127] ^ data[128] ^ data[129] ^ data[130] ^ data[131] ^ data[133] ^ data[134] ^ data[136] ^ data[137] ^ data[139] ^ data[141] ^ data[144] ^ data[145] ^ data[147] ^ data[148] ^ data[149] ^ data[150] ^ data[156] ^ data[157] ^ data[158] ^ data[159] ^ data[165] ^ data[166] ^ data[167] ^ data[168] ^ data[169] ^ data[171] ^ data[174] ^ data[175] ^ data[177] ^ data[179] ^ data[180] ^ data[181] ^ data[185] ^ data[188] ^ data[190] ^ data[192] ^ data[194] ^ data[195] ^ data[197] ^ data[199] ^ data[200] ^ data[201] ^ data[207] ^ data[209] ^ data[211] ^ data[212] ^ data[215] ^ data[218] ^ data[223] ^ data[224] ^ data[225] ^ data[228] ^ data[229] ^ data[231] ^ data[233] ^ data[234] ^ data[235] ^ data[238] ^ data[239] ^ data[240] ^ data[241] ^ data[244] ^ data[245] ^ data[246] ^ data[249] ^ data[250] ^ data[252] ;

assign temp_checkbits0[21] = checkbits[1] ^ checkbits[2] ^ checkbits[4] ^ checkbits[5] ^ checkbits[7] ^ checkbits[8] ^ checkbits[9] ^ checkbits[12] ^ checkbits[15] ^ checkbits[16] ^ checkbits[19] ^ checkbits[20] ^ checkbits[21] ^ checkbits[22] ^ checkbits[25] ^ checkbits[29] ^ checkbits[32] ^ checkbits[33] ^ data[0] ^ data[3] ^ data[5] ^ data[6] ^ data[8] ^ data[9] ^ data[10] ^ data[12] ^ data[14] ^ data[15] ^ data[17] ^ data[19] ^ data[21] ^ data[23] ^ data[24] ^ data[25] ^ data[29] ^ data[35] ^ data[37] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[44] ^ data[46] ^ data[47] ^ data[49] ^ data[52] ^ data[53] ^ data[54] ^ data[58] ^ data[60] ^ data[61] ^ data[63] ^ data[64] ^ data[67] ^ data[68] ^ data[70] ^ data[74] ^ data[75] ^ data[76] ^ data[77] ^ data[78] ^ data[79] ^ data[81] ^ data[85] ^ data[87] ^ data[88] ^ data[95] ^ data[100] ^ data[102] ^ data[104] ^ data[106] ^ data[108] ^ data[109] ^ data[112] ^ data[113] ^ data[116] ^ data[118] ^ data[119] ^ data[120] ^ data[121] ^ data[123] ^ data[124] ^ data[125] ^ data[128] ^ data[129] ^ data[130] ^ data[131] ^ data[132] ^ data[134] ^ data[135] ^ data[137] ^ data[138] ^ data[140] ^ data[142] ^ data[145] ^ data[146] ^ data[148] ^ data[149] ^ data[150] ^ data[151] ^ data[157] ^ data[158] ^ data[159] ^ data[160] ^ data[166] ^ data[167] ^ data[168] ^ data[169] ^ data[170] ^ data[172] ^ data[175] ^ data[176] ^ data[178] ^ data[180] ^ data[181] ^ data[182] ^ data[186] ^ data[189] ^ data[191] ^ data[193] ^ data[195] ^ data[196] ^ data[198] ^ data[200] ^ data[201] ^ data[202] ^ data[208] ^ data[210] ^ data[212] ^ data[213] ^ data[216] ^ data[219] ^ data[224] ^ data[225] ^ data[226] ^ data[229] ^ data[230] ^ data[232] ^ data[234] ^ data[235] ^ data[236] ^ data[239] ^ data[240] ^ data[241] ^ data[242] ^ data[245] ^ data[246] ^ data[247] ^ data[250] ^ data[251] ^ data[253] ;


assign temp_checkbits0[20] = checkbits[0] ^ checkbits[1] ^ checkbits[3] ^ checkbits[4] ^ checkbits[6] ^ checkbits[7] ^ checkbits[8] ^ checkbits[11] ^ checkbits[14] ^ checkbits[15] ^ checkbits[18] ^ checkbits[19] ^ checkbits[20] ^ checkbits[21] ^ checkbits[24] ^ checkbits[28] ^ checkbits[31] ^ checkbits[32] ^ data[1] ^ data[4] ^ data[6] ^ data[7] ^ data[9] ^ data[10] ^ data[11] ^ data[13] ^ data[15] ^ data[16] ^ data[18] ^ data[20] ^ data[22] ^ data[24] ^ data[25] ^ data[26] ^ data[30] ^ data[36] ^ data[38] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[45] ^ data[47] ^ data[48] ^ data[50] ^ data[53] ^ data[54] ^ data[55] ^ data[59] ^ data[61] ^ data[62] ^ data[64] ^ data[65] ^ data[68] ^ data[69] ^ data[71] ^ data[75] ^ data[76] ^ data[77] ^ data[78] ^ data[79] ^ data[80] ^ data[82] ^ data[86] ^ data[88] ^ data[89] ^ data[96] ^ data[101] ^ data[103] ^ data[105] ^ data[107] ^ data[109] ^ data[110] ^ data[113] ^ data[114] ^ data[117] ^ data[119] ^ data[120] ^ data[121] ^ data[122] ^ data[124] ^ data[125] ^ data[126] ^ data[129] ^ data[130] ^ data[131] ^ data[132] ^ data[133] ^ data[135] ^ data[136] ^ data[138] ^ data[139] ^ data[141] ^ data[143] ^ data[146] ^ data[147] ^ data[149] ^ data[150] ^ data[151] ^ data[152] ^ data[158] ^ data[159] ^ data[160] ^ data[161] ^ data[167] ^ data[168] ^ data[169] ^ data[170] ^ data[171] ^ data[173] ^ data[176] ^ data[177] ^ data[179] ^ data[181] ^ data[182] ^ data[183] ^ data[187] ^ data[190] ^ data[192] ^ data[194] ^ data[196] ^ data[197] ^ data[199] ^ data[201] ^ data[202] ^ data[203] ^ data[209] ^ data[211] ^ data[213] ^ data[214] ^ data[217] ^ data[220] ^ data[225] ^ data[226] ^ data[227] ^ data[230] ^ data[231] ^ data[233] ^ data[235] ^ data[236] ^ data[237] ^ data[240] ^ data[241] ^ data[242] ^ data[243] ^ data[246] ^ data[247] ^ data[248] ^ data[251] ^ data[252] ^ data[254] ;

assign temp_checkbits0[19] = checkbits[0] ^ checkbits[2] ^ checkbits[3] ^ checkbits[5] ^ checkbits[6] ^ checkbits[7] ^ checkbits[10] ^ checkbits[13] ^ checkbits[14] ^ checkbits[17] ^ checkbits[18] ^ checkbits[19] ^ checkbits[20] ^ checkbits[23] ^ checkbits[27] ^ checkbits[30] ^ checkbits[31] ^ data[0] ^ data[2] ^ data[5] ^ data[7] ^ data[8] ^ data[10] ^ data[11] ^ data[12] ^ data[14] ^ data[16] ^ data[17] ^ data[19] ^ data[21] ^ data[23] ^ data[25] ^ data[26] ^ data[27] ^ data[31] ^ data[37] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[46] ^ data[48] ^ data[49] ^ data[51] ^ data[54] ^ data[55] ^ data[56] ^ data[60] ^ data[62] ^ data[63] ^ data[65] ^ data[66] ^ data[69] ^ data[70] ^ data[72] ^ data[76] ^ data[77] ^ data[78] ^ data[79] ^ data[80] ^ data[81] ^ data[83] ^ data[87] ^ data[89] ^ data[90] ^ data[97] ^ data[102] ^ data[104] ^ data[106] ^ data[108] ^ data[110] ^ data[111] ^ data[114] ^ data[115] ^ data[118] ^ data[120] ^ data[121] ^ data[122] ^ data[123] ^ data[125] ^ data[126] ^ data[127] ^ data[130] ^ data[131] ^ data[132] ^ data[133] ^ data[134] ^ data[136] ^ data[137] ^ data[139] ^ data[140] ^ data[142] ^ data[144] ^ data[147] ^ data[148] ^ data[150] ^ data[151] ^ data[152] ^ data[153] ^ data[159] ^ data[160] ^ data[161] ^ data[162] ^ data[168] ^ data[169] ^ data[170] ^ data[171] ^ data[172] ^ data[174] ^ data[177] ^ data[178] ^ data[180] ^ data[182] ^ data[183] ^ data[184] ^ data[188] ^ data[191] ^ data[193] ^ data[195] ^ data[197] ^ data[198] ^ data[200] ^ data[202] ^ data[203] ^ data[204] ^ data[210] ^ data[212] ^ data[214] ^ data[215] ^ data[218] ^ data[221] ^ data[226] ^ data[227] ^ data[228] ^ data[231] ^ data[232] ^ data[234] ^ data[236] ^ data[237] ^ data[238] ^ data[241] ^ data[242] ^ data[243] ^ data[244] ^ data[247] ^ data[248] ^ data[249] ^ data[252] ^ data[253] ^ data[255] ;

assign temp_checkbits0[18] = checkbits[2] ^ checkbits[3] ^ checkbits[6] ^ checkbits[7] ^ checkbits[8] ^ checkbits[9] ^ checkbits[10] ^ checkbits[11] ^ checkbits[13] ^ checkbits[14] ^ checkbits[15] ^ checkbits[16] ^ checkbits[18] ^ checkbits[25] ^ checkbits[27] ^ checkbits[28] ^ checkbits[31] ^ checkbits[32] ^ data[0] ^ data[1] ^ data[2] ^ data[5] ^ data[6] ^ data[9] ^ data[10] ^ data[11] ^ data[19] ^ data[20] ^ data[21] ^ data[23] ^ data[24] ^ data[25] ^ data[26] ^ data[27] ^ data[28] ^ data[31] ^ data[32] ^ data[33] ^ data[35] ^ data[37] ^ data[40] ^ data[42] ^ data[44] ^ data[46] ^ data[47] ^ data[56] ^ data[59] ^ data[62] ^ data[67] ^ data[68] ^ data[69] ^ data[70] ^ data[71] ^ data[73] ^ data[78] ^ data[79] ^ data[80] ^ data[82] ^ data[84] ^ data[85] ^ data[86] ^ data[88] ^ data[90] ^ data[91] ^ data[93] ^ data[95] ^ data[97] ^ data[99] ^ data[100] ^ data[102] ^ data[104] ^ data[108] ^ data[109] ^ data[115] ^ data[116] ^ data[120] ^ data[121] ^ data[126] ^ data[128] ^ data[130] ^ data[131] ^ data[133] ^ data[136] ^ data[139] ^ data[140] ^ data[142] ^ data[145] ^ data[146] ^ data[149] ^ data[152] ^ data[155] ^ data[156] ^ data[157] ^ data[158] ^ data[160] ^ data[161] ^ data[162] ^ data[163] ^ data[166] ^ data[167] ^ data[168] ^ data[169] ^ data[173] ^ data[175] ^ data[176] ^ data[177] ^ data[179] ^ data[181] ^ data[182] ^ data[184] ^ data[185] ^ data[188] ^ data[189] ^ data[195] ^ data[197] ^ data[198] ^ data[201] ^ data[203] ^ data[205] ^ data[207] ^ data[210] ^ data[213] ^ data[215] ^ data[216] ^ data[218] ^ data[220] ^ data[223] ^ data[225] ^ data[226] ^ data[227] ^ data[228] ^ data[229] ^ data[237] ^ data[238] ^ data[241] ^ data[243] ^ data[246] ^ data[247] ^ data[248] ^ data[249] ^ data[250] ^ data[251] ^ data[252] ^ data[254] ;

assign temp_checkbits0[17] = checkbits[2] ^ checkbits[3] ^ checkbits[4] ^ checkbits[6] ^ checkbits[9] ^ checkbits[11] ^ checkbits[13] ^ checkbits[19] ^ checkbits[22] ^ checkbits[24] ^ checkbits[25] ^ checkbits[28] ^ checkbits[29] ^ checkbits[32] ^ data[1] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[11] ^ data[13] ^ data[15] ^ data[17] ^ data[18] ^ data[19] ^ data[20] ^ data[23] ^ data[24] ^ data[26] ^ data[27] ^ data[28] ^ data[29] ^ data[31] ^ data[32] ^ data[34] ^ data[35] ^ data[36] ^ data[37] ^ data[45] ^ data[46] ^ data[47] ^ data[48] ^ data[49] ^ data[50] ^ data[52] ^ data[55] ^ data[59] ^ data[60] ^ data[61] ^ data[62] ^ data[64] ^ data[66] ^ data[70] ^ data[71] ^ data[72] ^ data[74] ^ data[77] ^ data[79] ^ data[80] ^ data[83] ^ data[87] ^ data[89] ^ data[91] ^ data[92] ^ data[93] ^ data[94] ^ data[95] ^ data[96] ^ data[97] ^ data[99] ^ data[101] ^ data[102] ^ data[104] ^ data[107] ^ data[108] ^ data[109] ^ data[110] ^ data[111] ^ data[112] ^ data[116] ^ data[117] ^ data[119] ^ data[120] ^ data[121] ^ data[123] ^ data[124] ^ data[129] ^ data[130] ^ data[131] ^ data[135] ^ data[136] ^ data[138] ^ data[139] ^ data[140] ^ data[142] ^ data[147] ^ data[148] ^ data[150] ^ data[151] ^ data[154] ^ data[155] ^ data[159] ^ data[161] ^ data[162] ^ data[163] ^ data[164] ^ data[166] ^ data[169] ^ data[171] ^ data[172] ^ data[174] ^ data[180] ^ data[185] ^ data[186] ^ data[188] ^ data[189] ^ data[190] ^ data[192] ^ data[194] ^ data[195] ^ data[197] ^ data[198] ^ data[202] ^ data[206] ^ data[207] ^ data[208] ^ data[210] ^ data[214] ^ data[216] ^ data[217] ^ data[218] ^ data[220] ^ data[221] ^ data[222] ^ data[223] ^ data[224] ^ data[225] ^ data[227] ^ data[228] ^ data[229] ^ data[230] ^ data[232] ^ data[233] ^ data[235] ^ data[238] ^ data[241] ^ data[245] ^ data[246] ^ data[248] ^ data[249] ^ data[250] ^ data[255] ;

assign temp_checkbits0[16] = checkbits[2] ^ checkbits[4] ^ checkbits[7] ^ checkbits[11] ^ checkbits[14] ^ checkbits[15] ^ checkbits[17] ^ checkbits[18] ^ checkbits[19] ^ checkbits[21] ^ checkbits[22] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[29] ^ checkbits[30] ^ checkbits[32] ^ checkbits[35] ^ data[3] ^ data[5] ^ data[6] ^ data[7] ^ data[9] ^ data[10] ^ data[13] ^ data[14] ^ data[15] ^ data[16] ^ data[17] ^ data[20] ^ data[22] ^ data[23] ^ data[24] ^ data[27] ^ data[28] ^ data[29] ^ data[30] ^ data[31] ^ data[32] ^ data[36] ^ data[41] ^ data[43] ^ data[47] ^ data[48] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[56] ^ data[57] ^ data[59] ^ data[60] ^ data[64] ^ data[65] ^ data[66] ^ data[67] ^ data[68] ^ data[69] ^ data[71] ^ data[72] ^ data[73] ^ data[75] ^ data[77] ^ data[78] ^ data[80] ^ data[84] ^ data[85] ^ data[86] ^ data[88] ^ data[90] ^ data[92] ^ data[94] ^ data[96] ^ data[99] ^ data[104] ^ data[107] ^ data[109] ^ data[110] ^ data[113] ^ data[117] ^ data[118] ^ data[119] ^ data[121] ^ data[123] ^ data[125] ^ data[127] ^ data[131] ^ data[134] ^ data[135] ^ data[138] ^ data[140] ^ data[142] ^ data[146] ^ data[149] ^ data[152] ^ data[153] ^ data[154] ^ data[157] ^ data[158] ^ data[160] ^ data[162] ^ data[163] ^ data[164] ^ data[165] ^ data[166] ^ data[168] ^ data[171] ^ data[173] ^ data[175] ^ data[176] ^ data[177] ^ data[178] ^ data[181] ^ data[182] ^ data[183] ^ data[186] ^ data[187] ^ data[188] ^ data[189] ^ data[190] ^ data[191] ^ data[192] ^ data[193] ^ data[194] ^ data[197] ^ data[198] ^ data[203] ^ data[204] ^ data[208] ^ data[209] ^ data[210] ^ data[215] ^ data[217] ^ data[220] ^ data[221] ^ data[224] ^ data[228] ^ data[229] ^ data[230] ^ data[231] ^ data[232] ^ data[234] ^ data[235] ^ data[236] ^ data[241] ^ data[244] ^ data[245] ^ data[249] ^ data[250] ^ data[252] ^ data[253] ;

assign temp_checkbits0[15] = checkbits[1] ^ checkbits[3] ^ checkbits[6] ^ checkbits[10] ^ checkbits[13] ^ checkbits[14] ^ checkbits[16] ^ checkbits[17] ^ checkbits[18] ^ checkbits[20] ^ checkbits[21] ^ checkbits[22] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[28] ^ checkbits[29] ^ checkbits[31] ^ checkbits[34] ^ data[4] ^ data[6] ^ data[7] ^ data[8] ^ data[10] ^ data[11] ^ data[14] ^ data[15] ^ data[16] ^ data[17] ^ data[18] ^ data[21] ^ data[23] ^ data[24] ^ data[25] ^ data[28] ^ data[29] ^ data[30] ^ data[31] ^ data[32] ^ data[33] ^ data[37] ^ data[42] ^ data[44] ^ data[48] ^ data[49] ^ data[52] ^ data[53] ^ data[54] ^ data[56] ^ data[57] ^ data[58] ^ data[60] ^ data[61] ^ data[65] ^ data[66] ^ data[67] ^ data[68] ^ data[69] ^ data[70] ^ data[72] ^ data[73] ^ data[74] ^ data[76] ^ data[78] ^ data[79] ^ data[81] ^ data[85] ^ data[86] ^ data[87] ^ data[89] ^ data[91] ^ data[93] ^ data[95] ^ data[97] ^ data[100] ^ data[105] ^ data[108] ^ data[110] ^ data[111] ^ data[114] ^ data[118] ^ data[119] ^ data[120] ^ data[122] ^ data[124] ^ data[126] ^ data[128] ^ data[132] ^ data[135] ^ data[136] ^ data[139] ^ data[141] ^ data[143] ^ data[147] ^ data[150] ^ data[153] ^ data[154] ^ data[155] ^ data[158] ^ data[159] ^ data[161] ^ data[163] ^ data[164] ^ data[165] ^ data[166] ^ data[167] ^ data[169] ^ data[172] ^ data[174] ^ data[176] ^ data[177] ^ data[178] ^ data[179] ^ data[182] ^ data[183] ^ data[184] ^ data[187] ^ data[188] ^ data[189] ^ data[190] ^ data[191] ^ data[192] ^ data[193] ^ data[194] ^ data[195] ^ data[198] ^ data[199] ^ data[204] ^ data[205] ^ data[209] ^ data[210] ^ data[211] ^ data[216] ^ data[218] ^ data[221] ^ data[222] ^ data[225] ^ data[229] ^ data[230] ^ data[231] ^ data[232] ^ data[233] ^ data[235] ^ data[236] ^ data[237] ^ data[242] ^ data[245] ^ data[246] ^ data[250] ^ data[251] ^ data[253] ^ data[254] ;

assign temp_checkbits0[14] = checkbits[0] ^ checkbits[1] ^ checkbits[2] ^ checkbits[3] ^ checkbits[4] ^ checkbits[7] ^ checkbits[8] ^ checkbits[9] ^ checkbits[10] ^ checkbits[11] ^ checkbits[13] ^ checkbits[14] ^ checkbits[16] ^ checkbits[20] ^ checkbits[21] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[29] ^ checkbits[31] ^ checkbits[32] ^ checkbits[33] ^ checkbits[35] ^ data[2] ^ data[3] ^ data[7] ^ data[9] ^ data[10] ^ data[11] ^ data[13] ^ data[16] ^ data[21] ^ data[23] ^ data[24] ^ data[26] ^ data[29] ^ data[30] ^ data[32] ^ data[34] ^ data[35] ^ data[37] ^ data[41] ^ data[45] ^ data[46] ^ data[52] ^ data[53] ^ data[54] ^ data[58] ^ data[63] ^ data[64] ^ data[67] ^ data[70] ^ data[71] ^ data[73] ^ data[74] ^ data[75] ^ data[79] ^ data[80] ^ data[81] ^ data[82] ^ data[85] ^ data[87] ^ data[88] ^ data[90] ^ data[92] ^ data[93] ^ data[94] ^ data[95] ^ data[96] ^ data[97] ^ data[99] ^ data[100] ^ data[101] ^ data[102] ^ data[103] ^ data[104] ^ data[105] ^ data[106] ^ data[107] ^ data[108] ^ data[109] ^ data[115] ^ data[121] ^ data[122] ^ data[124] ^ data[125] ^ data[129] ^ data[130] ^ data[132] ^ data[133] ^ data[134] ^ data[135] ^ data[138] ^ data[139] ^ data[140] ^ data[141] ^ data[143] ^ data[144] ^ data[146] ^ data[153] ^ data[157] ^ data[158] ^ data[159] ^ data[160] ^ data[162] ^ data[164] ^ data[165] ^ data[171] ^ data[172] ^ data[173] ^ data[175] ^ data[176] ^ data[179] ^ data[180] ^ data[182] ^ data[184] ^ data[185] ^ data[189] ^ data[190] ^ data[191] ^ data[193] ^ data[197] ^ data[200] ^ data[204] ^ data[205] ^ data[206] ^ data[207] ^ data[212] ^ data[217] ^ data[218] ^ data[220] ^ data[225] ^ data[230] ^ data[231] ^ data[234] ^ data[235] ^ data[236] ^ data[237] ^ data[238] ^ data[239] ^ data[241] ^ data[242] ^ data[243] ^ data[244] ^ data[245] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[13] = checkbits[0] ^ checkbits[2] ^ checkbits[4] ^ checkbits[5] ^ checkbits[6] ^ checkbits[9] ^ checkbits[11] ^ checkbits[13] ^ checkbits[14] ^ checkbits[17] ^ checkbits[20] ^ checkbits[23] ^ checkbits[24] ^ checkbits[26] ^ checkbits[27] ^ checkbits[29] ^ checkbits[34] ^ data[0] ^ data[2] ^ data[4] ^ data[5] ^ data[11] ^ data[13] ^ data[14] ^ data[15] ^ data[18] ^ data[19] ^ data[21] ^ data[23] ^ data[24] ^ data[27] ^ data[30] ^ data[36] ^ data[37] ^ data[41] ^ data[42] ^ data[43] ^ data[47] ^ data[49] ^ data[50] ^ data[52] ^ data[53] ^ data[54] ^ data[57] ^ data[61] ^ data[62] ^ data[63] ^ data[65] ^ data[66] ^ data[69] ^ data[71] ^ data[72] ^ data[74] ^ data[75] ^ data[76] ^ data[77] ^ data[80] ^ data[82] ^ data[83] ^ data[85] ^ data[88] ^ data[89] ^ data[91] ^ data[94] ^ data[96] ^ data[99] ^ data[101] ^ data[106] ^ data[109] ^ data[110] ^ data[111] ^ data[112] ^ data[116] ^ data[119] ^ data[120] ^ data[124] ^ data[125] ^ data[126] ^ data[127] ^ data[131] ^ data[132] ^ data[133] ^ data[137] ^ data[138] ^ data[140] ^ data[143] ^ data[144] ^ data[145] ^ data[146] ^ data[147] ^ data[148] ^ data[151] ^ data[153] ^ data[155] ^ data[156] ^ data[157] ^ data[159] ^ data[160] ^ data[161] ^ data[163] ^ data[165] ^ data[167] ^ data[168] ^ data[170] ^ data[171] ^ data[173] ^ data[174] ^ data[178] ^ data[180] ^ data[181] ^ data[182] ^ data[185] ^ data[186] ^ data[188] ^ data[190] ^ data[191] ^ data[195] ^ data[196] ^ data[197] ^ data[198] ^ data[199] ^ data[201] ^ data[204] ^ data[205] ^ data[206] ^ data[208] ^ data[210] ^ data[211] ^ data[213] ^ data[220] ^ data[221] ^ data[222] ^ data[223] ^ data[225] ^ data[231] ^ data[233] ^ data[236] ^ data[237] ^ data[238] ^ data[240] ^ data[241] ^ data[243] ^ data[247] ^ data[251] ^ data[252] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[12] = checkbits[1] ^ checkbits[3] ^ checkbits[4] ^ checkbits[5] ^ checkbits[8] ^ checkbits[10] ^ checkbits[12] ^ checkbits[13] ^ checkbits[16] ^ checkbits[19] ^ checkbits[22] ^ checkbits[23] ^ checkbits[25] ^ checkbits[26] ^ checkbits[28] ^ checkbits[33] ^ data[0] ^ data[1] ^ data[3] ^ data[5] ^ data[6] ^ data[12] ^ data[14] ^ data[15] ^ data[16] ^ data[19] ^ data[20] ^ data[22] ^ data[24] ^ data[25] ^ data[28] ^ data[31] ^ data[37] ^ data[38] ^ data[42] ^ data[43] ^ data[44] ^ data[48] ^ data[50] ^ data[51] ^ data[53] ^ data[54] ^ data[55] ^ data[58] ^ data[62] ^ data[63] ^ data[64] ^ data[66] ^ data[67] ^ data[70] ^ data[72] ^ data[73] ^ data[75] ^ data[76] ^ data[77] ^ data[78] ^ data[81] ^ data[83] ^ data[84] ^ data[86] ^ data[89] ^ data[90] ^ data[92] ^ data[95] ^ data[97] ^ data[100] ^ data[102] ^ data[107] ^ data[110] ^ data[111] ^ data[112] ^ data[113] ^ data[117] ^ data[120] ^ data[121] ^ data[125] ^ data[126] ^ data[127] ^ data[128] ^ data[132] ^ data[133] ^ data[134] ^ data[138] ^ data[139] ^ data[141] ^ data[144] ^ data[145] ^ data[146] ^ data[147] ^ data[148] ^ data[149] ^ data[152] ^ data[154] ^ data[156] ^ data[157] ^ data[158] ^ data[160] ^ data[161] ^ data[162] ^ data[164] ^ data[166] ^ data[168] ^ data[169] ^ data[171] ^ data[172] ^ data[174] ^ data[175] ^ data[179] ^ data[181] ^ data[182] ^ data[183] ^ data[186] ^ data[187] ^ data[189] ^ data[191] ^ data[192] ^ data[196] ^ data[197] ^ data[198] ^ data[199] ^ data[200] ^ data[202] ^ data[205] ^ data[206] ^ data[207] ^ data[209] ^ data[211] ^ data[212] ^ data[214] ^ data[221] ^ data[222] ^ data[223] ^ data[224] ^ data[226] ^ data[232] ^ data[234] ^ data[237] ^ data[238] ^ data[239] ^ data[241] ^ data[242] ^ data[244] ^ data[248] ^ data[252] ^ data[253] ^ data[254] ^ data[255] ;

assign temp_checkbits0[11] = checkbits[0] ^ checkbits[1] ^ checkbits[2] ^ checkbits[5] ^ checkbits[8] ^ checkbits[9] ^ checkbits[10] ^ checkbits[14] ^ checkbits[17] ^ checkbits[18] ^ checkbits[19] ^ checkbits[21] ^ checkbits[24] ^ checkbits[26] ^ checkbits[28] ^ checkbits[29] ^ checkbits[30] ^ checkbits[31] ^ data[1] ^ data[3] ^ data[4] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[10] ^ data[12] ^ data[16] ^ data[18] ^ data[19] ^ data[20] ^ data[22] ^ data[26] ^ data[29] ^ data[31] ^ data[32] ^ data[33] ^ data[35] ^ data[37] ^ data[39] ^ data[41] ^ data[44] ^ data[45] ^ data[46] ^ data[50] ^ data[51] ^ data[54] ^ data[56] ^ data[57] ^ data[61] ^ data[62] ^ data[65] ^ data[66] ^ data[67] ^ data[69] ^ data[71] ^ data[73] ^ data[74] ^ data[76] ^ data[78] ^ data[79] ^ data[81] ^ data[82] ^ data[84] ^ data[86] ^ data[87] ^ data[90] ^ data[91] ^ data[95] ^ data[96] ^ data[97] ^ data[99] ^ data[100] ^ data[101] ^ data[102] ^ data[104] ^ data[105] ^ data[107] ^ data[113] ^ data[114] ^ data[118] ^ data[119] ^ data[120] ^ data[121] ^ data[123] ^ data[124] ^ data[126] ^ data[128] ^ data[129] ^ data[130] ^ data[132] ^ data[133] ^ data[136] ^ data[137] ^ data[138] ^ data[140] ^ data[141] ^ data[143] ^ data[145] ^ data[147] ^ data[149] ^ data[150] ^ data[151] ^ data[154] ^ data[156] ^ data[159] ^ data[161] ^ data[162] ^ data[163] ^ data[165] ^ data[166] ^ data[168] ^ data[169] ^ data[171] ^ data[173] ^ data[175] ^ data[177] ^ data[178] ^ data[180] ^ data[184] ^ data[187] ^ data[190] ^ data[193] ^ data[194] ^ data[195] ^ data[196] ^ data[198] ^ data[200] ^ data[201] ^ data[203] ^ data[204] ^ data[206] ^ data[208] ^ data[211] ^ data[212] ^ data[213] ^ data[215] ^ data[218] ^ data[219] ^ data[220] ^ data[224] ^ data[226] ^ data[227] ^ data[232] ^ data[238] ^ data[240] ^ data[241] ^ data[243] ^ data[244] ^ data[246] ^ data[247] ^ data[249] ^ data[251] ^ data[252] ^ data[254] ^ data[255] ;

assign temp_checkbits0[10] = checkbits[0] ^ checkbits[1] ^ checkbits[4] ^ checkbits[7] ^ checkbits[8] ^ checkbits[9] ^ checkbits[13] ^ checkbits[16] ^ checkbits[17] ^ checkbits[18] ^ checkbits[20] ^ checkbits[23] ^ checkbits[25] ^ checkbits[27] ^ checkbits[28] ^ checkbits[29] ^ checkbits[30] ^ checkbits[35] ^ data[0] ^ data[2] ^ data[4] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[9] ^ data[11] ^ data[13] ^ data[17] ^ data[19] ^ data[20] ^ data[21] ^ data[23] ^ data[27] ^ data[30] ^ data[32] ^ data[33] ^ data[34] ^ data[36] ^ data[38] ^ data[40] ^ data[42] ^ data[45] ^ data[46] ^ data[47] ^ data[51] ^ data[52] ^ data[55] ^ data[57] ^ data[58] ^ data[62] ^ data[63] ^ data[66] ^ data[67] ^ data[68] ^ data[70] ^ data[72] ^ data[74] ^ data[75] ^ data[77] ^ data[79] ^ data[80] ^ data[82] ^ data[83] ^ data[85] ^ data[87] ^ data[88] ^ data[91] ^ data[92] ^ data[96] ^ data[97] ^ data[98] ^ data[100] ^ data[101] ^ data[102] ^ data[103] ^ data[105] ^ data[106] ^ data[108] ^ data[114] ^ data[115] ^ data[119] ^ data[120] ^ data[121] ^ data[122] ^ data[124] ^ data[125] ^ data[127] ^ data[129] ^ data[130] ^ data[131] ^ data[133] ^ data[134] ^ data[137] ^ data[138] ^ data[139] ^ data[141] ^ data[142] ^ data[144] ^ data[146] ^ data[148] ^ data[150] ^ data[151] ^ data[152] ^ data[155] ^ data[157] ^ data[160] ^ data[162] ^ data[163] ^ data[164] ^ data[166] ^ data[167] ^ data[169] ^ data[170] ^ data[172] ^ data[174] ^ data[176] ^ data[178] ^ data[179] ^ data[181] ^ data[185] ^ data[188] ^ data[191] ^ data[194] ^ data[195] ^ data[196] ^ data[197] ^ data[199] ^ data[201] ^ data[202] ^ data[204] ^ data[205] ^ data[207] ^ data[209] ^ data[212] ^ data[213] ^ data[214] ^ data[216] ^ data[219] ^ data[220] ^ data[221] ^ data[225] ^ data[227] ^ data[228] ^ data[233] ^ data[239] ^ data[241] ^ data[242] ^ data[244] ^ data[245] ^ data[247] ^ data[248] ^ data[250] ^ data[252] ^ data[253] ^ data[255] ;

assign temp_checkbits0[9] = checkbits[0] ^ checkbits[3] ^ checkbits[6] ^ checkbits[7] ^ checkbits[8] ^ checkbits[12] ^ checkbits[15] ^ checkbits[16] ^ checkbits[17] ^ checkbits[19] ^ checkbits[22] ^ checkbits[24] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[29] ^ checkbits[34] ^ data[0] ^ data[1] ^ data[3] ^ data[5] ^ data[6] ^ data[7] ^ data[8] ^ data[9] ^ data[10] ^ data[12] ^ data[14] ^ data[18] ^ data[20] ^ data[21] ^ data[22] ^ data[24] ^ data[28] ^ data[31] ^ data[33] ^ data[34] ^ data[35] ^ data[37] ^ data[39] ^ data[41] ^ data[43] ^ data[46] ^ data[47] ^ data[48] ^ data[52] ^ data[53] ^ data[56] ^ data[58] ^ data[59] ^ data[63] ^ data[64] ^ data[67] ^ data[68] ^ data[69] ^ data[71] ^ data[73] ^ data[75] ^ data[76] ^ data[78] ^ data[80] ^ data[81] ^ data[83] ^ data[84] ^ data[86] ^ data[88] ^ data[89] ^ data[92] ^ data[93] ^ data[97] ^ data[98] ^ data[99] ^ data[101] ^ data[102] ^ data[103] ^ data[104] ^ data[106] ^ data[107] ^ data[109] ^ data[115] ^ data[116] ^ data[120] ^ data[121] ^ data[122] ^ data[123] ^ data[125] ^ data[126] ^ data[128] ^ data[130] ^ data[131] ^ data[132] ^ data[134] ^ data[135] ^ data[138] ^ data[139] ^ data[140] ^ data[142] ^ data[143] ^ data[145] ^ data[147] ^ data[149] ^ data[151] ^ data[152] ^ data[153] ^ data[156] ^ data[158] ^ data[161] ^ data[163] ^ data[164] ^ data[165] ^ data[167] ^ data[168] ^ data[170] ^ data[171] ^ data[173] ^ data[175] ^ data[177] ^ data[179] ^ data[180] ^ data[182] ^ data[186] ^ data[189] ^ data[192] ^ data[195] ^ data[196] ^ data[197] ^ data[198] ^ data[200] ^ data[202] ^ data[203] ^ data[205] ^ data[206] ^ data[208] ^ data[210] ^ data[213] ^ data[214] ^ data[215] ^ data[217] ^ data[220] ^ data[221] ^ data[222] ^ data[226] ^ data[228] ^ data[229] ^ data[234] ^ data[240] ^ data[242] ^ data[243] ^ data[245] ^ data[246] ^ data[248] ^ data[249] ^ data[251] ^ data[253] ^ data[254] ;

assign temp_checkbits0[8] = checkbits[2] ^ checkbits[5] ^ checkbits[6] ^ checkbits[7] ^ checkbits[11] ^ checkbits[14] ^ checkbits[15] ^ checkbits[16] ^ checkbits[18] ^ checkbits[21] ^ checkbits[23] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[33] ^ data[0] ^ data[1] ^ data[2] ^ data[4] ^ data[6] ^ data[7] ^ data[8] ^ data[9] ^ data[10] ^ data[11] ^ data[13] ^ data[15] ^ data[19] ^ data[21] ^ data[22] ^ data[23] ^ data[25] ^ data[29] ^ data[32] ^ data[34] ^ data[35] ^ data[36] ^ data[38] ^ data[40] ^ data[42] ^ data[44] ^ data[47] ^ data[48] ^ data[49] ^ data[53] ^ data[54] ^ data[57] ^ data[59] ^ data[60] ^ data[64] ^ data[65] ^ data[68] ^ data[69] ^ data[70] ^ data[72] ^ data[74] ^ data[76] ^ data[77] ^ data[79] ^ data[81] ^ data[82] ^ data[84] ^ data[85] ^ data[87] ^ data[89] ^ data[90] ^ data[93] ^ data[94] ^ data[98] ^ data[99] ^ data[100] ^ data[102] ^ data[103] ^ data[104] ^ data[105] ^ data[107] ^ data[108] ^ data[110] ^ data[116] ^ data[117] ^ data[121] ^ data[122] ^ data[123] ^ data[124] ^ data[126] ^ data[127] ^ data[129] ^ data[131] ^ data[132] ^ data[133] ^ data[135] ^ data[136] ^ data[139] ^ data[140] ^ data[141] ^ data[143] ^ data[144] ^ data[146] ^ data[148] ^ data[150] ^ data[152] ^ data[153] ^ data[154] ^ data[157] ^ data[159] ^ data[162] ^ data[164] ^ data[165] ^ data[166] ^ data[168] ^ data[169] ^ data[171] ^ data[172] ^ data[174] ^ data[176] ^ data[178] ^ data[180] ^ data[181] ^ data[183] ^ data[187] ^ data[190] ^ data[193] ^ data[196] ^ data[197] ^ data[198] ^ data[199] ^ data[201] ^ data[203] ^ data[204] ^ data[206] ^ data[207] ^ data[209] ^ data[211] ^ data[214] ^ data[215] ^ data[216] ^ data[218] ^ data[221] ^ data[222] ^ data[223] ^ data[227] ^ data[229] ^ data[230] ^ data[235] ^ data[241] ^ data[243] ^ data[244] ^ data[246] ^ data[247] ^ data[249] ^ data[250] ^ data[252] ^ data[254] ^ data[255] ;

assign temp_checkbits0[7] = checkbits[1] ^ checkbits[4] ^ checkbits[5] ^ checkbits[6] ^ checkbits[10] ^ checkbits[13] ^ checkbits[14] ^ checkbits[15] ^ checkbits[17] ^ checkbits[20] ^ checkbits[22] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[32] ^ data[1] ^ data[2] ^ data[3] ^ data[5] ^ data[7] ^ data[8] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[14] ^ data[16] ^ data[20] ^ data[22] ^ data[23] ^ data[24] ^ data[26] ^ data[30] ^ data[33] ^ data[35] ^ data[36] ^ data[37] ^ data[39] ^ data[41] ^ data[43] ^ data[45] ^ data[48] ^ data[49] ^ data[50] ^ data[54] ^ data[55] ^ data[58] ^ data[60] ^ data[61] ^ data[65] ^ data[66] ^ data[69] ^ data[70] ^ data[71] ^ data[73] ^ data[75] ^ data[77] ^ data[78] ^ data[80] ^ data[82] ^ data[83] ^ data[85] ^ data[86] ^ data[88] ^ data[90] ^ data[91] ^ data[94] ^ data[95] ^ data[99] ^ data[100] ^ data[101] ^ data[103] ^ data[104] ^ data[105] ^ data[106] ^ data[108] ^ data[109] ^ data[111] ^ data[117] ^ data[118] ^ data[122] ^ data[123] ^ data[124] ^ data[125] ^ data[127] ^ data[128] ^ data[130] ^ data[132] ^ data[133] ^ data[134] ^ data[136] ^ data[137] ^ data[140] ^ data[141] ^ data[142] ^ data[144] ^ data[145] ^ data[147] ^ data[149] ^ data[151] ^ data[153] ^ data[154] ^ data[155] ^ data[158] ^ data[160] ^ data[163] ^ data[165] ^ data[166] ^ data[167] ^ data[169] ^ data[170] ^ data[172] ^ data[173] ^ data[175] ^ data[177] ^ data[179] ^ data[181] ^ data[182] ^ data[184] ^ data[188] ^ data[191] ^ data[194] ^ data[197] ^ data[198] ^ data[199] ^ data[200] ^ data[202] ^ data[204] ^ data[205] ^ data[207] ^ data[208] ^ data[210] ^ data[212] ^ data[215] ^ data[216] ^ data[217] ^ data[219] ^ data[222] ^ data[223] ^ data[224] ^ data[228] ^ data[230] ^ data[231] ^ data[236] ^ data[242] ^ data[244] ^ data[245] ^ data[247] ^ data[248] ^ data[250] ^ data[251] ^ data[253] ^ data[255] ;

assign temp_checkbits0[6] = checkbits[0] ^ checkbits[3] ^ checkbits[4] ^ checkbits[5] ^ checkbits[9] ^ checkbits[12] ^ checkbits[13] ^ checkbits[14] ^ checkbits[16] ^ checkbits[19] ^ checkbits[21] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[31] ^ checkbits[35] ^ data[2] ^ data[3] ^ data[4] ^ data[6] ^ data[8] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[15] ^ data[17] ^ data[21] ^ data[23] ^ data[24] ^ data[25] ^ data[27] ^ data[31] ^ data[34] ^ data[36] ^ data[37] ^ data[38] ^ data[40] ^ data[42] ^ data[44] ^ data[46] ^ data[49] ^ data[50] ^ data[51] ^ data[55] ^ data[56] ^ data[59] ^ data[61] ^ data[62] ^ data[66] ^ data[67] ^ data[70] ^ data[71] ^ data[72] ^ data[74] ^ data[76] ^ data[78] ^ data[79] ^ data[81] ^ data[83] ^ data[84] ^ data[86] ^ data[87] ^ data[89] ^ data[91] ^ data[92] ^ data[95] ^ data[96] ^ data[100] ^ data[101] ^ data[102] ^ data[104] ^ data[105] ^ data[106] ^ data[107] ^ data[109] ^ data[110] ^ data[112] ^ data[118] ^ data[119] ^ data[123] ^ data[124] ^ data[125] ^ data[126] ^ data[128] ^ data[129] ^ data[131] ^ data[133] ^ data[134] ^ data[135] ^ data[137] ^ data[138] ^ data[141] ^ data[142] ^ data[143] ^ data[145] ^ data[146] ^ data[148] ^ data[150] ^ data[152] ^ data[154] ^ data[155] ^ data[156] ^ data[159] ^ data[161] ^ data[164] ^ data[166] ^ data[167] ^ data[168] ^ data[170] ^ data[171] ^ data[173] ^ data[174] ^ data[176] ^ data[178] ^ data[180] ^ data[182] ^ data[183] ^ data[185] ^ data[189] ^ data[192] ^ data[195] ^ data[198] ^ data[199] ^ data[200] ^ data[201] ^ data[203] ^ data[205] ^ data[206] ^ data[208] ^ data[209] ^ data[211] ^ data[213] ^ data[216] ^ data[217] ^ data[218] ^ data[220] ^ data[223] ^ data[224] ^ data[225] ^ data[229] ^ data[231] ^ data[232] ^ data[237] ^ data[243] ^ data[245] ^ data[246] ^ data[248] ^ data[249] ^ data[251] ^ data[252] ^ data[254] ;

assign temp_checkbits0[5] = checkbits[2] ^ checkbits[3] ^ checkbits[4] ^ checkbits[8] ^ checkbits[11] ^ checkbits[12] ^ checkbits[13] ^ checkbits[15] ^ checkbits[18] ^ checkbits[20] ^ checkbits[22] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[30] ^ checkbits[34] ^ checkbits[35] ^ data[0] ^ data[3] ^ data[4] ^ data[5] ^ data[7] ^ data[9] ^ data[10] ^ data[11] ^ data[12] ^ data[13] ^ data[14] ^ data[16] ^ data[18] ^ data[22] ^ data[24] ^ data[25] ^ data[26] ^ data[28] ^ data[32] ^ data[35] ^ data[37] ^ data[38] ^ data[39] ^ data[41] ^ data[43] ^ data[45] ^ data[47] ^ data[50] ^ data[51] ^ data[52] ^ data[56] ^ data[57] ^ data[60] ^ data[62] ^ data[63] ^ data[67] ^ data[68] ^ data[71] ^ data[72] ^ data[73] ^ data[75] ^ data[77] ^ data[79] ^ data[80] ^ data[82] ^ data[84] ^ data[85] ^ data[87] ^ data[88] ^ data[90] ^ data[92] ^ data[93] ^ data[96] ^ data[97] ^ data[101] ^ data[102] ^ data[103] ^ data[105] ^ data[106] ^ data[107] ^ data[108] ^ data[110] ^ data[111] ^ data[113] ^ data[119] ^ data[120] ^ data[124] ^ data[125] ^ data[126] ^ data[127] ^ data[129] ^ data[130] ^ data[132] ^ data[134] ^ data[135] ^ data[136] ^ data[138] ^ data[139] ^ data[142] ^ data[143] ^ data[144] ^ data[146] ^ data[147] ^ data[149] ^ data[151] ^ data[153] ^ data[155] ^ data[156] ^ data[157] ^ data[160] ^ data[162] ^ data[165] ^ data[167] ^ data[168] ^ data[169] ^ data[171] ^ data[172] ^ data[174] ^ data[175] ^ data[177] ^ data[179] ^ data[181] ^ data[183] ^ data[184] ^ data[186] ^ data[190] ^ data[193] ^ data[196] ^ data[199] ^ data[200] ^ data[201] ^ data[202] ^ data[204] ^ data[206] ^ data[207] ^ data[209] ^ data[210] ^ data[212] ^ data[214] ^ data[217] ^ data[218] ^ data[219] ^ data[221] ^ data[224] ^ data[225] ^ data[226] ^ data[230] ^ data[232] ^ data[233] ^ data[238] ^ data[244] ^ data[246] ^ data[247] ^ data[249] ^ data[250] ^ data[252] ^ data[253] ^ data[255] ;

assign temp_checkbits0[4] = checkbits[2] ^ checkbits[4] ^ checkbits[5] ^ checkbits[8] ^ checkbits[15] ^ checkbits[21] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[30] ^ checkbits[31] ^ checkbits[32] ^ checkbits[33] ^ checkbits[34] ^ checkbits[35] ^ data[1] ^ data[2] ^ data[3] ^ data[4] ^ data[6] ^ data[11] ^ data[14] ^ data[18] ^ data[21] ^ data[22] ^ data[26] ^ data[27] ^ data[29] ^ data[31] ^ data[35] ^ data[36] ^ data[37] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[48] ^ data[49] ^ data[50] ^ data[51] ^ data[53] ^ data[55] ^ data[58] ^ data[59] ^ data[62] ^ data[66] ^ data[72] ^ data[73] ^ data[74] ^ data[76] ^ data[77] ^ data[78] ^ data[80] ^ data[83] ^ data[88] ^ data[89] ^ data[91] ^ data[94] ^ data[95] ^ data[99] ^ data[100] ^ data[105] ^ data[106] ^ data[109] ^ data[114] ^ data[119] ^ data[121] ^ data[122] ^ data[123] ^ data[124] ^ data[125] ^ data[126] ^ data[128] ^ data[131] ^ data[132] ^ data[133] ^ data[134] ^ data[138] ^ data[140] ^ data[141] ^ data[142] ^ data[144] ^ data[145] ^ data[146] ^ data[147] ^ data[150] ^ data[151] ^ data[152] ^ data[153] ^ data[155] ^ data[161] ^ data[163] ^ data[167] ^ data[169] ^ data[171] ^ data[173] ^ data[175] ^ data[177] ^ data[180] ^ data[183] ^ data[184] ^ data[185] ^ data[187] ^ data[188] ^ data[191] ^ data[192] ^ data[195] ^ data[196] ^ data[199] ^ data[200] ^ data[201] ^ data[202] ^ data[203] ^ data[204] ^ data[205] ^ data[208] ^ data[213] ^ data[215] ^ data[223] ^ data[227] ^ data[231] ^ data[232] ^ data[234] ^ data[235] ^ data[241] ^ data[242] ^ data[244] ^ data[246] ^ data[248] ^ data[250] ^ data[252] ^ data[254] ;

assign temp_checkbits0[3] = checkbits[1] ^ checkbits[3] ^ checkbits[4] ^ checkbits[7] ^ checkbits[14] ^ checkbits[20] ^ checkbits[22] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[27] ^ checkbits[29] ^ checkbits[30] ^ checkbits[31] ^ checkbits[32] ^ checkbits[33] ^ checkbits[34] ^ data[2] ^ data[3] ^ data[4] ^ data[5] ^ data[7] ^ data[12] ^ data[15] ^ data[19] ^ data[22] ^ data[23] ^ data[27] ^ data[28] ^ data[30] ^ data[32] ^ data[36] ^ data[37] ^ data[38] ^ data[40] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[49] ^ data[50] ^ data[51] ^ data[52] ^ data[54] ^ data[56] ^ data[59] ^ data[60] ^ data[63] ^ data[67] ^ data[73] ^ data[74] ^ data[75] ^ data[77] ^ data[78] ^ data[79] ^ data[81] ^ data[84] ^ data[89] ^ data[90] ^ data[92] ^ data[95] ^ data[96] ^ data[100] ^ data[101] ^ data[106] ^ data[107] ^ data[110] ^ data[115] ^ data[120] ^ data[122] ^ data[123] ^ data[124] ^ data[125] ^ data[126] ^ data[127] ^ data[129] ^ data[132] ^ data[133] ^ data[134] ^ data[135] ^ data[139] ^ data[141] ^ data[142] ^ data[143] ^ data[145] ^ data[146] ^ data[147] ^ data[148] ^ data[151] ^ data[152] ^ data[153] ^ data[154] ^ data[156] ^ data[162] ^ data[164] ^ data[168] ^ data[170] ^ data[172] ^ data[174] ^ data[176] ^ data[178] ^ data[181] ^ data[184] ^ data[185] ^ data[186] ^ data[188] ^ data[189] ^ data[192] ^ data[193] ^ data[196] ^ data[197] ^ data[200] ^ data[201] ^ data[202] ^ data[203] ^ data[204] ^ data[205] ^ data[206] ^ data[209] ^ data[214] ^ data[216] ^ data[224] ^ data[228] ^ data[232] ^ data[233] ^ data[235] ^ data[236] ^ data[242] ^ data[243] ^ data[245] ^ data[247] ^ data[249] ^ data[251] ^ data[253] ^ data[255] ;

assign temp_checkbits0[2] = checkbits[0] ^ checkbits[2] ^ checkbits[3] ^ checkbits[6] ^ checkbits[13] ^ checkbits[19] ^ checkbits[21] ^ checkbits[22] ^ checkbits[23] ^ checkbits[24] ^ checkbits[25] ^ checkbits[26] ^ checkbits[28] ^ checkbits[29] ^ checkbits[30] ^ checkbits[31] ^ checkbits[32] ^ checkbits[33] ^ checkbits[35] ^ data[3] ^ data[4] ^ data[5] ^ data[6] ^ data[8] ^ data[13] ^ data[16] ^ data[20] ^ data[23] ^ data[24] ^ data[28] ^ data[29] ^ data[31] ^ data[33] ^ data[37] ^ data[38] ^ data[39] ^ data[41] ^ data[42] ^ data[43] ^ data[44] ^ data[45] ^ data[46] ^ data[50] ^ data[51] ^ data[52] ^ data[53] ^ data[55] ^ data[57] ^ data[60] ^ data[61] ^ data[64] ^ data[68] ^ data[74] ^ data[75] ^ data[76] ^ data[78] ^ data[79] ^ data[80] ^ data[82] ^ data[85] ^ data[90] ^ data[91] ^ data[93] ^ data[96] ^ data[97] ^ data[101] ^ data[102] ^ data[107] ^ data[108] ^ data[111] ^ data[116] ^ data[121] ^ data[123] ^ data[124] ^ data[125] ^ data[126] ^ data[127] ^ data[128] ^ data[130] ^ data[133] ^ data[134] ^ data[135] ^ data[136] ^ data[140] ^ data[142] ^ data[143] ^ data[144] ^ data[146] ^ data[147] ^ data[148] ^ data[149] ^ data[152] ^ data[153] ^ data[154] ^ data[155] ^ data[157] ^ data[163] ^ data[165] ^ data[169] ^ data[171] ^ data[173] ^ data[175] ^ data[177] ^ data[179] ^ data[182] ^ data[185] ^ data[186] ^ data[187] ^ data[189] ^ data[190] ^ data[193] ^ data[194] ^ data[197] ^ data[198] ^ data[201] ^ data[202] ^ data[203] ^ data[204] ^ data[205] ^ data[206] ^ data[207] ^ data[210] ^ data[215] ^ data[217] ^ data[225] ^ data[229] ^ data[233] ^ data[234] ^ data[236] ^ data[237] ^ data[243] ^ data[244] ^ data[246] ^ data[248] ^ data[250] ^ data[252] ^ data[254] ;

assign temp_checkbits0[1] = checkbits[2] ^ checkbits[3] ^ checkbits[4] ^ checkbits[7] ^ checkbits[8] ^ checkbits[10] ^ checkbits[11] ^ checkbits[14] ^ checkbits[15] ^ checkbits[17] ^ checkbits[18] ^ checkbits[19] ^ checkbits[20] ^ checkbits[21] ^ checkbits[23] ^ checkbits[24] ^ checkbits[26] ^ checkbits[34] ^ data[0] ^ data[2] ^ data[3] ^ data[4] ^ data[6] ^ data[7] ^ data[8] ^ data[9] ^ data[10] ^ data[12] ^ data[13] ^ data[14] ^ data[15] ^ data[18] ^ data[19] ^ data[22] ^ data[23] ^ data[24] ^ data[29] ^ data[30] ^ data[31] ^ data[32] ^ data[33] ^ data[34] ^ data[35] ^ data[37] ^ data[39] ^ data[40] ^ data[41] ^ data[42] ^ data[44] ^ data[45] ^ data[47] ^ data[49] ^ data[50] ^ data[51] ^ data[53] ^ data[54] ^ data[55] ^ data[56] ^ data[57] ^ data[58] ^ data[59] ^ data[63] ^ data[64] ^ data[65] ^ data[66] ^ data[68] ^ data[75] ^ data[76] ^ data[79] ^ data[80] ^ data[83] ^ data[85] ^ data[91] ^ data[92] ^ data[93] ^ data[94] ^ data[95] ^ data[99] ^ data[100] ^ data[104] ^ data[105] ^ data[107] ^ data[109] ^ data[111] ^ data[117] ^ data[119] ^ data[120] ^ data[123] ^ data[125] ^ data[126] ^ data[128] ^ data[129] ^ data[130] ^ data[131] ^ data[132] ^ data[138] ^ data[139] ^ data[142] ^ data[144] ^ data[145] ^ data[146] ^ data[147] ^ data[149] ^ data[150] ^ data[151] ^ data[157] ^ data[164] ^ data[167] ^ data[168] ^ data[171] ^ data[174] ^ data[177] ^ data[180] ^ data[182] ^ data[186] ^ data[187] ^ data[190] ^ data[191] ^ data[192] ^ data[196] ^ data[197] ^ data[198] ^ data[202] ^ data[203] ^ data[205] ^ data[206] ^ data[208] ^ data[210] ^ data[216] ^ data[219] ^ data[220] ^ data[222] ^ data[223] ^ data[225] ^ data[230] ^ data[232] ^ data[233] ^ data[234] ^ data[237] ^ data[238] ^ data[239] ^ data[241] ^ data[242] ^ data[246] ^ data[249] ^ data[252] ^ data[255] ;

assign temp_checkbits0[0] = checkbits[2] ^ checkbits[4] ^ checkbits[5] ^ checkbits[6] ^ checkbits[8] ^ checkbits[9] ^ checkbits[11] ^ checkbits[12] ^ checkbits[13] ^ checkbits[15] ^ checkbits[16] ^ checkbits[18] ^ checkbits[20] ^ checkbits[23] ^ checkbits[26] ^ checkbits[27] ^ checkbits[28] ^ checkbits[29] ^ checkbits[30] ^ checkbits[31] ^ checkbits[32] ^ checkbits[33] ^ data[1] ^ data[2] ^ data[4] ^ data[7] ^ data[9] ^ data[11] ^ data[12] ^ data[14] ^ data[16] ^ data[17] ^ data[18] ^ data[20] ^ data[21] ^ data[22] ^ data[24] ^ data[30] ^ data[32] ^ data[34] ^ data[36] ^ data[37] ^ data[40] ^ data[42] ^ data[45] ^ data[48] ^ data[49] ^ data[51] ^ data[54] ^ data[56] ^ data[58] ^ data[60] ^ data[61] ^ data[62] ^ data[63] ^ data[65] ^ data[67] ^ data[68] ^ data[76] ^ data[80] ^ data[84] ^ data[85] ^ data[92] ^ data[94] ^ data[96] ^ data[97] ^ data[98] ^ data[99] ^ data[101] ^ data[102] ^ data[103] ^ data[104] ^ data[106] ^ data[107] ^ data[110] ^ data[111] ^ data[118] ^ data[119] ^ data[121] ^ data[122] ^ data[123] ^ data[126] ^ data[129] ^ data[131] ^ data[133] ^ data[134] ^ data[135] ^ data[136] ^ data[137] ^ data[138] ^ data[140] ^ data[141] ^ data[142] ^ data[145] ^ data[147] ^ data[150] ^ data[152] ^ data[153] ^ data[154] ^ data[155] ^ data[156] ^ data[157] ^ data[165] ^ data[166] ^ data[167] ^ data[169] ^ data[170] ^ data[171] ^ data[175] ^ data[176] ^ data[177] ^ data[181] ^ data[182] ^ data[187] ^ data[191] ^ data[193] ^ data[194] ^ data[195] ^ data[196] ^ data[198] ^ data[203] ^ data[206] ^ data[209] ^ data[210] ^ data[217] ^ data[218] ^ data[219] ^ data[221] ^ data[222] ^ data[224] ^ data[225] ^ data[231] ^ data[232] ^ data[234] ^ data[238] ^ data[240] ^ data[241] ^ data[243] ^ data[244] ^ data[245] ^ data[246] ^ data[250] ^ data[251] ^ data[252] ;




assign temp_checkbits1[35] =   data[257] ^ data[258] ^ data[259] ^ data[262] ^ data[263] ^ data[265] ^ data[267] ^ data[268] ^ data[272] ^ data[273] ^ data[274] ^ data[276] ^ data[277] ^ data[278] ^ data[282] ^ data[285] ^ data[287] ^ data[288] ^ data[291] ^ data[293] ^ data[294] ^ data[298] ^ data[299] ^ data[300] ^ data[302] ^ data[303] ^ data[304] ^ data[305] ^ data[306] ^ data[308] ^ data[310] ^ data[311] ^ data[312] ^ data[315] ^ data[320] ^ data[321] ^ data[323] ^ data[324] ^ data[326] ^ data[327] ^ data[329] ^ data[330] ^ data[335] ^ data[338] ^ data[342] ^ data[346] ^ data[349] ^ data[351] ^ data[355] ^ data[356] ^ data[357] ^ data[358] ^ data[364] ^ data[369] ^ data[372] ^ data[373] ^ data[374] ^ data[376] ^ data[378] ^ data[379] ^ data[380] ^ data[381] ^ data[382] ^ data[383] ^ data[385] ^ data[386] ^ data[387] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[393] ^ data[394] ^ data[395] ^ data[396] ^ data[398] ^ data[399] ^ data[405] ^ data[410] ^ data[411] ^ data[412] ^ data[414] ^ data[418] ^ data[420] ^ data[423] ^ data[424] ^ data[426] ^ data[433] ^ data[435] ^ data[436] ^ data[442] ^ data[444] ^ data[446] ^ data[447] ^ data[450] ^ data[452] ^ data[453] ^ data[454] ^ data[455] ^ data[460] ^ data[461] ^ data[462] ^ data[466] ^ data[468] ^ data[471] ^ data[472] ^ data[474] ^ data[476];

assign temp_checkbits1[34] =   data[258] ^ data[259] ^ data[260] ^ data[263] ^ data[264] ^ data[266] ^ data[268] ^ data[269] ^ data[273] ^ data[274] ^ data[275] ^ data[277] ^ data[278] ^ data[279] ^ data[283] ^ data[286] ^ data[288] ^ data[289] ^ data[292] ^ data[294] ^ data[295] ^ data[299] ^ data[300] ^ data[301] ^ data[303] ^ data[304] ^ data[305] ^ data[306] ^ data[307] ^ data[309] ^ data[311] ^ data[312] ^ data[313] ^ data[316] ^ data[321] ^ data[322] ^ data[324] ^ data[325] ^ data[327] ^ data[328] ^ data[330] ^ data[331] ^ data[336] ^ data[339] ^ data[343] ^ data[347] ^ data[350] ^ data[352] ^ data[356] ^ data[357] ^ data[358] ^ data[359] ^ data[365] ^ data[370] ^ data[373] ^ data[374] ^ data[375] ^ data[377] ^ data[379] ^ data[380] ^ data[381] ^ data[382] ^ data[383] ^ data[384] ^ data[386] ^ data[387] ^ data[388] ^ data[390] ^ data[391] ^ data[392] ^ data[393] ^ data[394] ^ data[395] ^ data[396] ^ data[397] ^ data[399] ^ data[400] ^ data[406] ^ data[411] ^ data[412] ^ data[413] ^ data[415] ^ data[419] ^ data[421] ^ data[424] ^ data[425] ^ data[427] ^ data[434] ^ data[436] ^ data[437] ^ data[443] ^ data[445] ^ data[447] ^ data[448] ^ data[451] ^ data[453] ^ data[454] ^ data[455] ^ data[456] ^ data[461] ^ data[462] ^ data[463] ^ data[467] ^ data[469] ^ data[472] ^ data[473] ^ data[475] ^ data[477];

assign temp_checkbits1[33] =   data[257] ^ data[258] ^ data[260] ^ data[261] ^ data[262] ^ data[263] ^ data[264] ^ data[268] ^ data[269] ^ data[270] ^ data[272] ^ data[273] ^ data[275] ^ data[277] ^ data[279] ^ data[280] ^ data[282] ^ data[284] ^ data[285] ^ data[288] ^ data[289] ^ data[290] ^ data[291] ^ data[294] ^ data[295] ^ data[296] ^ data[298] ^ data[299] ^ data[301] ^ data[303] ^ data[307] ^ data[311] ^ data[313] ^ data[314] ^ data[315] ^ data[317] ^ data[320] ^ data[321] ^ data[322] ^ data[324] ^ data[325] ^ data[327] ^ data[328] ^ data[330] ^ data[331] ^ data[332] ^ data[335] ^ data[337] ^ data[338] ^ data[340] ^ data[342] ^ data[344] ^ data[346] ^ data[348] ^ data[349] ^ data[353] ^ data[355] ^ data[356] ^ data[359] ^ data[360] ^ data[364] ^ data[366] ^ data[369] ^ data[371] ^ data[372] ^ data[373] ^ data[375] ^ data[379] ^ data[384] ^ data[386] ^ data[388] ^ data[390] ^ data[397] ^ data[399] ^ data[400] ^ data[401] ^ data[405] ^ data[407] ^ data[410] ^ data[411] ^ data[413] ^ data[416] ^ data[418] ^ data[422] ^ data[423] ^ data[424] ^ data[425] ^ data[428] ^ data[433] ^ data[436] ^ data[437] ^ data[438] ^ data[442] ^ data[447] ^ data[448] ^ data[449] ^ data[450] ^ data[453] ^ data[456] ^ data[457] ^ data[460] ^ data[461] ^ data[463] ^ data[464] ^ data[466] ^ data[470] ^ data[471] ^ data[472] ^ data[473] ^ data[478];

assign temp_checkbits1[32] =   data[256] ^ data[258] ^ data[259] ^ data[261] ^ data[262] ^ data[263] ^ data[264] ^ data[265] ^ data[269] ^ data[270] ^ data[271] ^ data[273] ^ data[274] ^ data[276] ^ data[278] ^ data[280] ^ data[281] ^ data[283] ^ data[285] ^ data[286] ^ data[289] ^ data[290] ^ data[291] ^ data[292] ^ data[295] ^ data[296] ^ data[297] ^ data[299] ^ data[300] ^ data[302] ^ data[304] ^ data[308] ^ data[312] ^ data[314] ^ data[315] ^ data[316] ^ data[318] ^ data[321] ^ data[322] ^ data[323] ^ data[325] ^ data[326] ^ data[328] ^ data[329] ^ data[331] ^ data[332] ^ data[333] ^ data[336] ^ data[338] ^ data[339] ^ data[341] ^ data[343] ^ data[345] ^ data[347] ^ data[349] ^ data[350] ^ data[354] ^ data[356] ^ data[357] ^ data[360] ^ data[361] ^ data[365] ^ data[367] ^ data[370] ^ data[372] ^ data[373] ^ data[374] ^ data[376] ^ data[380] ^ data[385] ^ data[387] ^ data[389] ^ data[391] ^ data[398] ^ data[400] ^ data[401] ^ data[402] ^ data[406] ^ data[408] ^ data[411] ^ data[412] ^ data[414] ^ data[417] ^ data[419] ^ data[423] ^ data[424] ^ data[425] ^ data[426] ^ data[429] ^ data[434] ^ data[437] ^ data[438] ^ data[439] ^ data[443] ^ data[448] ^ data[449] ^ data[450] ^ data[451] ^ data[454] ^ data[457] ^ data[458] ^ data[461] ^ data[462] ^ data[464] ^ data[465] ^ data[467] ^ data[471] ^ data[472] ^ data[473] ^ data[474] ^ data[479];

assign temp_checkbits1[31] =   data[256] ^ data[257] ^ data[259] ^ data[260] ^ data[262] ^ data[263] ^ data[264] ^ data[265] ^ data[266] ^ data[270] ^ data[271] ^ data[272] ^ data[274] ^ data[275] ^ data[277] ^ data[279] ^ data[281] ^ data[282] ^ data[284] ^ data[286] ^ data[287] ^ data[290] ^ data[291] ^ data[292] ^ data[293] ^ data[296] ^ data[297] ^ data[298] ^ data[300] ^ data[301] ^ data[303] ^ data[305] ^ data[309] ^ data[313] ^ data[315] ^ data[316] ^ data[317] ^ data[319] ^ data[322] ^ data[323] ^ data[324] ^ data[326] ^ data[327] ^ data[329] ^ data[330] ^ data[332] ^ data[333] ^ data[334] ^ data[337] ^ data[339] ^ data[340] ^ data[342] ^ data[344] ^ data[346] ^ data[348] ^ data[350] ^ data[351] ^ data[355] ^ data[357] ^ data[358] ^ data[361] ^ data[362] ^ data[366] ^ data[368] ^ data[371] ^ data[373] ^ data[374] ^ data[375] ^ data[377] ^ data[381] ^ data[386] ^ data[388] ^ data[390] ^ data[392] ^ data[399] ^ data[401] ^ data[402] ^ data[403] ^ data[407] ^ data[409] ^ data[412] ^ data[413] ^ data[415] ^ data[418] ^ data[420] ^ data[424] ^ data[425] ^ data[426] ^ data[427] ^ data[430] ^ data[435] ^ data[438] ^ data[439] ^ data[440] ^ data[444] ^ data[449] ^ data[450] ^ data[451] ^ data[452] ^ data[455] ^ data[458] ^ data[459] ^ data[462] ^ data[463] ^ data[465] ^ data[466] ^ data[468] ^ data[472] ^ data[473] ^ data[474] ^ data[475] ^ data[480];

assign temp_checkbits1[30] =   data[259] ^ data[260] ^ data[261] ^ data[262] ^ data[264] ^ data[266] ^ data[268] ^ data[271] ^ data[274] ^ data[275] ^ data[277] ^ data[280] ^ data[283] ^ data[292] ^ data[297] ^ data[300] ^ data[301] ^ data[303] ^ data[305] ^ data[308] ^ data[311] ^ data[312] ^ data[314] ^ data[315] ^ data[316] ^ data[317] ^ data[318] ^ data[321] ^ data[325] ^ data[326] ^ data[328] ^ data[329] ^ data[331] ^ data[333] ^ data[334] ^ data[340] ^ data[341] ^ data[342] ^ data[343] ^ data[345] ^ data[346] ^ data[347] ^ data[352] ^ data[355] ^ data[357] ^ data[359] ^ data[362] ^ data[363] ^ data[364] ^ data[367] ^ data[373] ^ data[375] ^ data[379] ^ data[380] ^ data[381] ^ data[383] ^ data[385] ^ data[386] ^ data[390] ^ data[392] ^ data[394] ^ data[395] ^ data[396] ^ data[398] ^ data[399] ^ data[400] ^ data[402] ^ data[403] ^ data[404] ^ data[405] ^ data[408] ^ data[411] ^ data[412] ^ data[413] ^ data[416] ^ data[418] ^ data[419] ^ data[420] ^ data[421] ^ data[423] ^ data[424] ^ data[425] ^ data[427] ^ data[428] ^ data[431] ^ data[433] ^ data[435] ^ data[439] ^ data[440] ^ data[441] ^ data[442] ^ data[444] ^ data[445] ^ data[446] ^ data[447] ^ data[451] ^ data[454] ^ data[455] ^ data[456] ^ data[459] ^ data[461] ^ data[462] ^ data[463] ^ data[464] ^ data[467] ^ data[468] ^ data[469] ^ data[471] ^ data[472] ^ data[473] ^ data[475] ^ data[481];

assign temp_checkbits1[29] =   data[256] ^ data[257] ^ data[258] ^ data[259] ^ data[260] ^ data[261] ^ data[268] ^ data[269] ^ data[273] ^ data[274] ^ data[275] ^ data[277] ^ data[281] ^ data[282] ^ data[284] ^ data[285] ^ data[287] ^ data[288] ^ data[291] ^ data[294] ^ data[299] ^ data[300] ^ data[301] ^ data[303] ^ data[305] ^ data[308] ^ data[309] ^ data[310] ^ data[311] ^ data[313] ^ data[316] ^ data[317] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[332] ^ data[334] ^ data[338] ^ data[341] ^ data[343] ^ data[344] ^ data[347] ^ data[348] ^ data[349] ^ data[351] ^ data[353] ^ data[355] ^ data[357] ^ data[360] ^ data[363] ^ data[365] ^ data[368] ^ data[369] ^ data[372] ^ data[373] ^ data[378] ^ data[379] ^ data[383] ^ data[384] ^ data[385] ^ data[389] ^ data[390] ^ data[392] ^ data[394] ^ data[397] ^ data[398] ^ data[400] ^ data[401] ^ data[403] ^ data[404] ^ data[406] ^ data[409] ^ data[410] ^ data[411] ^ data[413] ^ data[417] ^ data[418] ^ data[419] ^ data[421] ^ data[422] ^ data[423] ^ data[425] ^ data[428] ^ data[429] ^ data[432] ^ data[433] ^ data[434] ^ data[435] ^ data[440] ^ data[441] ^ data[443] ^ data[444] ^ data[445] ^ data[448] ^ data[450] ^ data[453] ^ data[454] ^ data[456] ^ data[457] ^ data[461] ^ data[463] ^ data[464] ^ data[465] ^ data[466] ^ data[469] ^ data[470] ^ data[471] ^ data[473] ^ data[482];

assign temp_checkbits1[28] =   data[256] ^ data[257] ^ data[258] ^ data[259] ^ data[260] ^ data[261] ^ data[262] ^ data[269] ^ data[270] ^ data[274] ^ data[275] ^ data[276] ^ data[278] ^ data[282] ^ data[283] ^ data[285] ^ data[286] ^ data[288] ^ data[289] ^ data[292] ^ data[295] ^ data[300] ^ data[301] ^ data[302] ^ data[304] ^ data[306] ^ data[309] ^ data[310] ^ data[311] ^ data[312] ^ data[314] ^ data[317] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[333] ^ data[335] ^ data[339] ^ data[342] ^ data[344] ^ data[345] ^ data[348] ^ data[349] ^ data[350] ^ data[352] ^ data[354] ^ data[356] ^ data[358] ^ data[361] ^ data[364] ^ data[366] ^ data[369] ^ data[370] ^ data[373] ^ data[374] ^ data[379] ^ data[380] ^ data[384] ^ data[385] ^ data[386] ^ data[390] ^ data[391] ^ data[393] ^ data[395] ^ data[398] ^ data[399] ^ data[401] ^ data[402] ^ data[404] ^ data[405] ^ data[407] ^ data[410] ^ data[411] ^ data[412] ^ data[414] ^ data[418] ^ data[419] ^ data[420] ^ data[422] ^ data[423] ^ data[424] ^ data[426] ^ data[429] ^ data[430] ^ data[433] ^ data[434] ^ data[435] ^ data[436] ^ data[441] ^ data[442] ^ data[444] ^ data[445] ^ data[446] ^ data[449] ^ data[451] ^ data[454] ^ data[455] ^ data[457] ^ data[458] ^ data[462] ^ data[464] ^ data[465] ^ data[466] ^ data[467] ^ data[470] ^ data[471] ^ data[472] ^ data[474] ^ data[483];

assign temp_checkbits1[27] =   data[256] ^ data[257] ^ data[258] ^ data[259] ^ data[260] ^ data[261] ^ data[262] ^ data[263] ^ data[270] ^ data[271] ^ data[275] ^ data[276] ^ data[277] ^ data[279] ^ data[283] ^ data[284] ^ data[286] ^ data[287] ^ data[289] ^ data[290] ^ data[293] ^ data[296] ^ data[301] ^ data[302] ^ data[303] ^ data[305] ^ data[307] ^ data[310] ^ data[311] ^ data[312] ^ data[313] ^ data[315] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[334] ^ data[336] ^ data[340] ^ data[343] ^ data[345] ^ data[346] ^ data[349] ^ data[350] ^ data[351] ^ data[353] ^ data[355] ^ data[357] ^ data[359] ^ data[362] ^ data[365] ^ data[367] ^ data[370] ^ data[371] ^ data[374] ^ data[375] ^ data[380] ^ data[381] ^ data[385] ^ data[386] ^ data[387] ^ data[391] ^ data[392] ^ data[394] ^ data[396] ^ data[399] ^ data[400] ^ data[402] ^ data[403] ^ data[405] ^ data[406] ^ data[408] ^ data[411] ^ data[412] ^ data[413] ^ data[415] ^ data[419] ^ data[420] ^ data[421] ^ data[423] ^ data[424] ^ data[425] ^ data[427] ^ data[430] ^ data[431] ^ data[434] ^ data[435] ^ data[436] ^ data[437] ^ data[442] ^ data[443] ^ data[445] ^ data[446] ^ data[447] ^ data[450] ^ data[452] ^ data[455] ^ data[456] ^ data[458] ^ data[459] ^ data[463] ^ data[465] ^ data[466] ^ data[467] ^ data[468] ^ data[471] ^ data[472] ^ data[473] ^ data[475] ^ data[484];

assign temp_checkbits1[26] =   data[256] ^ data[260] ^ data[261] ^ data[264] ^ data[265] ^ data[267] ^ data[268] ^ data[271] ^ data[273] ^ data[274] ^ data[280] ^ data[282] ^ data[284] ^ data[290] ^ data[293] ^ data[297] ^ data[298] ^ data[299] ^ data[300] ^ data[305] ^ data[310] ^ data[313] ^ data[314] ^ data[315] ^ data[316] ^ data[319] ^ data[322] ^ data[325] ^ data[329] ^ data[330] ^ data[337] ^ data[338] ^ data[341] ^ data[342] ^ data[344] ^ data[347] ^ data[349] ^ data[350] ^ data[352] ^ data[354] ^ data[355] ^ data[357] ^ data[360] ^ data[363] ^ data[364] ^ data[366] ^ data[368] ^ data[369] ^ data[371] ^ data[373] ^ data[374] ^ data[375] ^ data[378] ^ data[379] ^ data[380] ^ data[383] ^ data[385] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[394] ^ data[396] ^ data[397] ^ data[398] ^ data[399] ^ data[400] ^ data[401] ^ data[403] ^ data[404] ^ data[405] ^ data[406] ^ data[407] ^ data[409] ^ data[410] ^ data[411] ^ data[413] ^ data[416] ^ data[418] ^ data[421] ^ data[422] ^ data[423] ^ data[425] ^ data[428] ^ data[431] ^ data[432] ^ data[433] ^ data[437] ^ data[438] ^ data[442] ^ data[443] ^ data[448] ^ data[450] ^ data[451] ^ data[452] ^ data[454] ^ data[455] ^ data[456] ^ data[457] ^ data[459] ^ data[461] ^ data[462] ^ data[464] ^ data[467] ^ data[469] ^ data[471] ^ data[473] ^ data[485];

assign temp_checkbits1[25] =   data[256] ^ data[257] ^ data[261] ^ data[262] ^ data[265] ^ data[266] ^ data[268] ^ data[269] ^ data[272] ^ data[274] ^ data[275] ^ data[281] ^ data[283] ^ data[285] ^ data[291] ^ data[294] ^ data[298] ^ data[299] ^ data[300] ^ data[301] ^ data[306] ^ data[311] ^ data[314] ^ data[315] ^ data[316] ^ data[317] ^ data[320] ^ data[323] ^ data[326] ^ data[330] ^ data[331] ^ data[338] ^ data[339] ^ data[342] ^ data[343] ^ data[345] ^ data[348] ^ data[350] ^ data[351] ^ data[353] ^ data[355] ^ data[356] ^ data[358] ^ data[361] ^ data[364] ^ data[365] ^ data[367] ^ data[369] ^ data[370] ^ data[372] ^ data[374] ^ data[375] ^ data[376] ^ data[379] ^ data[380] ^ data[381] ^ data[384] ^ data[386] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[395] ^ data[397] ^ data[398] ^ data[399] ^ data[400] ^ data[401] ^ data[402] ^ data[404] ^ data[405] ^ data[406] ^ data[407] ^ data[408] ^ data[410] ^ data[411] ^ data[412] ^ data[414] ^ data[417] ^ data[419] ^ data[422] ^ data[423] ^ data[424] ^ data[426] ^ data[429] ^ data[432] ^ data[433] ^ data[434] ^ data[438] ^ data[439] ^ data[443] ^ data[444] ^ data[449] ^ data[451] ^ data[452] ^ data[453] ^ data[455] ^ data[456] ^ data[457] ^ data[458] ^ data[460] ^ data[462] ^ data[463] ^ data[465] ^ data[468] ^ data[470] ^ data[472] ^ data[474] ^ data[486];

assign temp_checkbits1[24] =   data[256] ^ data[257] ^ data[258] ^ data[262] ^ data[263] ^ data[266] ^ data[267] ^ data[269] ^ data[270] ^ data[273] ^ data[275] ^ data[276] ^ data[282] ^ data[284] ^ data[286] ^ data[292] ^ data[295] ^ data[299] ^ data[300] ^ data[301] ^ data[302] ^ data[307] ^ data[312] ^ data[315] ^ data[316] ^ data[317] ^ data[318] ^ data[321] ^ data[324] ^ data[327] ^ data[331] ^ data[332] ^ data[339] ^ data[340] ^ data[343] ^ data[344] ^ data[346] ^ data[349] ^ data[351] ^ data[352] ^ data[354] ^ data[356] ^ data[357] ^ data[359] ^ data[362] ^ data[365] ^ data[366] ^ data[368] ^ data[370] ^ data[371] ^ data[373] ^ data[375] ^ data[376] ^ data[377] ^ data[380] ^ data[381] ^ data[382] ^ data[385] ^ data[387] ^ data[390] ^ data[391] ^ data[392] ^ data[393] ^ data[396] ^ data[398] ^ data[399] ^ data[400] ^ data[401] ^ data[402] ^ data[403] ^ data[405] ^ data[406] ^ data[407] ^ data[408] ^ data[409] ^ data[411] ^ data[412] ^ data[413] ^ data[415] ^ data[418] ^ data[420] ^ data[423] ^ data[424] ^ data[425] ^ data[427] ^ data[430] ^ data[433] ^ data[434] ^ data[435] ^ data[439] ^ data[440] ^ data[444] ^ data[445] ^ data[450] ^ data[452] ^ data[453] ^ data[454] ^ data[456] ^ data[457] ^ data[458] ^ data[459] ^ data[461] ^ data[463] ^ data[464] ^ data[466] ^ data[469] ^ data[471] ^ data[473] ^ data[475] ^ data[487];

assign temp_checkbits1[23] =   data[256] ^ data[262] ^ data[264] ^ data[265] ^ data[270] ^ data[271] ^ data[272] ^ data[273] ^ data[278] ^ data[282] ^ data[283] ^ data[288] ^ data[291] ^ data[294] ^ data[296] ^ data[298] ^ data[299] ^ data[301] ^ data[304] ^ data[305] ^ data[306] ^ data[310] ^ data[311] ^ data[312] ^ data[313] ^ data[315] ^ data[316] ^ data[317] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[332] ^ data[333] ^ data[335] ^ data[338] ^ data[340] ^ data[341] ^ data[342] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[349] ^ data[350] ^ data[351] ^ data[352] ^ data[353] ^ data[356] ^ data[360] ^ data[363] ^ data[364] ^ data[366] ^ data[367] ^ data[371] ^ data[373] ^ data[377] ^ data[379] ^ data[380] ^ data[385] ^ data[387] ^ data[388] ^ data[389] ^ data[390] ^ data[395] ^ data[396] ^ data[397] ^ data[398] ^ data[400] ^ data[401] ^ data[402] ^ data[403] ^ data[404] ^ data[405] ^ data[406] ^ data[407] ^ data[408] ^ data[409] ^ data[411] ^ data[413] ^ data[416] ^ data[418] ^ data[419] ^ data[420] ^ data[421] ^ data[423] ^ data[425] ^ data[428] ^ data[431] ^ data[433] ^ data[434] ^ data[440] ^ data[441] ^ data[442] ^ data[444] ^ data[445] ^ data[447] ^ data[450] ^ data[451] ^ data[452] ^ data[457] ^ data[458] ^ data[459] ^ data[461] ^ data[464] ^ data[465] ^ data[466] ^ data[467] ^ data[468] ^ data[470] ^ data[471] ^ data[488];

assign temp_checkbits1[22] =   data[257] ^ data[263] ^ data[265] ^ data[266] ^ data[271] ^ data[272] ^ data[273] ^ data[274] ^ data[279] ^ data[283] ^ data[284] ^ data[289] ^ data[292] ^ data[295] ^ data[297] ^ data[299] ^ data[300] ^ data[302] ^ data[305] ^ data[306] ^ data[307] ^ data[311] ^ data[312] ^ data[313] ^ data[314] ^ data[316] ^ data[317] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[331] ^ data[333] ^ data[334] ^ data[336] ^ data[339] ^ data[341] ^ data[342] ^ data[343] ^ data[345] ^ data[346] ^ data[347] ^ data[348] ^ data[350] ^ data[351] ^ data[352] ^ data[353] ^ data[354] ^ data[357] ^ data[361] ^ data[364] ^ data[365] ^ data[367] ^ data[368] ^ data[372] ^ data[374] ^ data[378] ^ data[380] ^ data[381] ^ data[386] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[396] ^ data[397] ^ data[398] ^ data[399] ^ data[401] ^ data[402] ^ data[403] ^ data[404] ^ data[405] ^ data[406] ^ data[407] ^ data[408] ^ data[409] ^ data[410] ^ data[412] ^ data[414] ^ data[417] ^ data[419] ^ data[420] ^ data[421] ^ data[422] ^ data[424] ^ data[426] ^ data[429] ^ data[432] ^ data[434] ^ data[435] ^ data[441] ^ data[442] ^ data[443] ^ data[445] ^ data[446] ^ data[448] ^ data[451] ^ data[452] ^ data[453] ^ data[458] ^ data[459] ^ data[460] ^ data[462] ^ data[465] ^ data[466] ^ data[467] ^ data[468] ^ data[469] ^ data[471] ^ data[472] ^ data[489];

assign temp_checkbits1[21] =   data[258] ^ data[264] ^ data[266] ^ data[267] ^ data[272] ^ data[273] ^ data[274] ^ data[275] ^ data[280] ^ data[284] ^ data[285] ^ data[290] ^ data[293] ^ data[296] ^ data[298] ^ data[300] ^ data[301] ^ data[303] ^ data[306] ^ data[307] ^ data[308] ^ data[312] ^ data[313] ^ data[314] ^ data[315] ^ data[317] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[331] ^ data[332] ^ data[334] ^ data[335] ^ data[337] ^ data[340] ^ data[342] ^ data[343] ^ data[344] ^ data[346] ^ data[347] ^ data[348] ^ data[349] ^ data[351] ^ data[352] ^ data[353] ^ data[354] ^ data[355] ^ data[358] ^ data[362] ^ data[365] ^ data[366] ^ data[368] ^ data[369] ^ data[373] ^ data[375] ^ data[379] ^ data[381] ^ data[382] ^ data[387] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[397] ^ data[398] ^ data[399] ^ data[400] ^ data[402] ^ data[403] ^ data[404] ^ data[405] ^ data[406] ^ data[407] ^ data[408] ^ data[409] ^ data[410] ^ data[411] ^ data[413] ^ data[415] ^ data[418] ^ data[420] ^ data[421] ^ data[422] ^ data[423] ^ data[425] ^ data[427] ^ data[430] ^ data[433] ^ data[435] ^ data[436] ^ data[442] ^ data[443] ^ data[444] ^ data[446] ^ data[447] ^ data[449] ^ data[452] ^ data[453] ^ data[454] ^ data[459] ^ data[460] ^ data[461] ^ data[463] ^ data[466] ^ data[467] ^ data[468] ^ data[469] ^ data[470] ^ data[472] ^ data[473] ^ data[490];

assign temp_checkbits1[20] =   data[259] ^ data[265] ^ data[267] ^ data[268] ^ data[273] ^ data[274] ^ data[275] ^ data[276] ^ data[281] ^ data[285] ^ data[286] ^ data[291] ^ data[294] ^ data[297] ^ data[299] ^ data[301] ^ data[302] ^ data[304] ^ data[307] ^ data[308] ^ data[309] ^ data[313] ^ data[314] ^ data[315] ^ data[316] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[331] ^ data[332] ^ data[333] ^ data[335] ^ data[336] ^ data[338] ^ data[341] ^ data[343] ^ data[344] ^ data[345] ^ data[347] ^ data[348] ^ data[349] ^ data[350] ^ data[352] ^ data[353] ^ data[354] ^ data[355] ^ data[356] ^ data[359] ^ data[363] ^ data[366] ^ data[367] ^ data[369] ^ data[370] ^ data[374] ^ data[376] ^ data[380] ^ data[382] ^ data[383] ^ data[388] ^ data[390] ^ data[391] ^ data[392] ^ data[393] ^ data[398] ^ data[399] ^ data[400] ^ data[401] ^ data[403] ^ data[404] ^ data[405] ^ data[406] ^ data[407] ^ data[408] ^ data[409] ^ data[410] ^ data[411] ^ data[412] ^ data[414] ^ data[416] ^ data[419] ^ data[421] ^ data[422] ^ data[423] ^ data[424] ^ data[426] ^ data[428] ^ data[431] ^ data[434] ^ data[436] ^ data[437] ^ data[443] ^ data[444] ^ data[445] ^ data[447] ^ data[448] ^ data[450] ^ data[453] ^ data[454] ^ data[455] ^ data[460] ^ data[461] ^ data[462] ^ data[464] ^ data[467] ^ data[468] ^ data[469] ^ data[470] ^ data[471] ^ data[473] ^ data[474] ^ data[491];

assign temp_checkbits1[19] =   data[260] ^ data[266] ^ data[268] ^ data[269] ^ data[274] ^ data[275] ^ data[276] ^ data[277] ^ data[282] ^ data[286] ^ data[287] ^ data[292] ^ data[295] ^ data[298] ^ data[300] ^ data[302] ^ data[303] ^ data[305] ^ data[308] ^ data[309] ^ data[310] ^ data[314] ^ data[315] ^ data[316] ^ data[317] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[331] ^ data[332] ^ data[333] ^ data[334] ^ data[336] ^ data[337] ^ data[339] ^ data[342] ^ data[344] ^ data[345] ^ data[346] ^ data[348] ^ data[349] ^ data[350] ^ data[351] ^ data[353] ^ data[354] ^ data[355] ^ data[356] ^ data[357] ^ data[360] ^ data[364] ^ data[367] ^ data[368] ^ data[370] ^ data[371] ^ data[375] ^ data[377] ^ data[381] ^ data[383] ^ data[384] ^ data[389] ^ data[391] ^ data[392] ^ data[393] ^ data[394] ^ data[399] ^ data[400] ^ data[401] ^ data[402] ^ data[404] ^ data[405] ^ data[406] ^ data[407] ^ data[408] ^ data[409] ^ data[410] ^ data[411] ^ data[412] ^ data[413] ^ data[415] ^ data[417] ^ data[420] ^ data[422] ^ data[423] ^ data[424] ^ data[425] ^ data[427] ^ data[429] ^ data[432] ^ data[435] ^ data[437] ^ data[438] ^ data[444] ^ data[445] ^ data[446] ^ data[448] ^ data[449] ^ data[451] ^ data[454] ^ data[455] ^ data[456] ^ data[461] ^ data[462] ^ data[463] ^ data[465] ^ data[468] ^ data[469] ^ data[470] ^ data[471] ^ data[472] ^ data[474] ^ data[475] ^ data[492];

assign temp_checkbits1[18] =   data[256] ^ data[257] ^ data[258] ^ data[259] ^ data[261] ^ data[262] ^ data[263] ^ data[265] ^ data[268] ^ data[269] ^ data[270] ^ data[272] ^ data[273] ^ data[274] ^ data[275] ^ data[282] ^ data[283] ^ data[285] ^ data[291] ^ data[294] ^ data[296] ^ data[298] ^ data[300] ^ data[301] ^ data[302] ^ data[305] ^ data[308] ^ data[309] ^ data[312] ^ data[316] ^ data[317] ^ data[318] ^ data[322] ^ data[325] ^ data[328] ^ data[331] ^ data[332] ^ data[333] ^ data[334] ^ data[337] ^ data[340] ^ data[342] ^ data[343] ^ data[345] ^ data[347] ^ data[350] ^ data[352] ^ data[354] ^ data[361] ^ data[364] ^ data[365] ^ data[368] ^ data[371] ^ data[373] ^ data[374] ^ data[379] ^ data[380] ^ data[381] ^ data[383] ^ data[384] ^ data[386] ^ data[387] ^ data[389] ^ data[391] ^ data[396] ^ data[398] ^ data[399] ^ data[400] ^ data[401] ^ data[402] ^ data[403] ^ data[406] ^ data[407] ^ data[408] ^ data[409] ^ data[413] ^ data[416] ^ data[420] ^ data[421] ^ data[425] ^ data[428] ^ data[430] ^ data[435] ^ data[438] ^ data[439] ^ data[442] ^ data[444] ^ data[445] ^ data[449] ^ data[453] ^ data[454] ^ data[456] ^ data[457] ^ data[460] ^ data[461] ^ data[463] ^ data[464] ^ data[468] ^ data[469] ^ data[470] ^ data[473] ^ data[474] ^ data[475] ^ data[493];

assign temp_checkbits1[17] =   data[260] ^ data[264] ^ data[265] ^ data[266] ^ data[267] ^ data[268] ^ data[269] ^ data[270] ^ data[271] ^ data[272] ^ data[275] ^ data[277] ^ data[278] ^ data[282] ^ data[283] ^ data[284] ^ data[285] ^ data[286] ^ data[287] ^ data[288] ^ data[291] ^ data[292] ^ data[293] ^ data[294] ^ data[295] ^ data[297] ^ data[298] ^ data[300] ^ data[301] ^ data[304] ^ data[305] ^ data[308] ^ data[309] ^ data[311] ^ data[312] ^ data[313] ^ data[315] ^ data[317] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[324] ^ data[327] ^ data[330] ^ data[332] ^ data[333] ^ data[334] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[348] ^ data[349] ^ data[353] ^ data[356] ^ data[357] ^ data[358] ^ data[362] ^ data[364] ^ data[365] ^ data[366] ^ data[373] ^ data[375] ^ data[376] ^ data[378] ^ data[379] ^ data[383] ^ data[384] ^ data[386] ^ data[388] ^ data[389] ^ data[391] ^ data[393] ^ data[394] ^ data[395] ^ data[396] ^ data[397] ^ data[398] ^ data[400] ^ data[401] ^ data[402] ^ data[403] ^ data[404] ^ data[405] ^ data[407] ^ data[408] ^ data[409] ^ data[411] ^ data[412] ^ data[417] ^ data[418] ^ data[420] ^ data[421] ^ data[422] ^ data[423] ^ data[424] ^ data[429] ^ data[431] ^ data[433] ^ data[435] ^ data[439] ^ data[440] ^ data[442] ^ data[443] ^ data[444] ^ data[445] ^ data[447] ^ data[452] ^ data[453] ^ data[457] ^ data[458] ^ data[460] ^ data[464] ^ data[465] ^ data[466] ^ data[468] ^ data[469] ^ data[470] ^ data[472] ^ data[475] ^ data[494];

assign temp_checkbits1[16] =   data[256] ^ data[257] ^ data[258] ^ data[259] ^ data[261] ^ data[262] ^ data[263] ^ data[266] ^ data[269] ^ data[270] ^ data[271] ^ data[274] ^ data[277] ^ data[279] ^ data[282] ^ data[283] ^ data[284] ^ data[286] ^ data[289] ^ data[291] ^ data[292] ^ data[295] ^ data[296] ^ data[300] ^ data[301] ^ data[303] ^ data[304] ^ data[308] ^ data[309] ^ data[311] ^ data[313] ^ data[314] ^ data[315] ^ data[316] ^ data[318] ^ data[319] ^ data[322] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[331] ^ data[333] ^ data[334] ^ data[338] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[350] ^ data[351] ^ data[354] ^ data[355] ^ data[356] ^ data[359] ^ data[363] ^ data[364] ^ data[365] ^ data[366] ^ data[367] ^ data[369] ^ data[372] ^ data[373] ^ data[377] ^ data[378] ^ data[381] ^ data[382] ^ data[383] ^ data[384] ^ data[386] ^ data[391] ^ data[393] ^ data[397] ^ data[401] ^ data[402] ^ data[403] ^ data[404] ^ data[406] ^ data[408] ^ data[409] ^ data[411] ^ data[413] ^ data[414] ^ data[419] ^ data[420] ^ data[421] ^ data[422] ^ data[425] ^ data[426] ^ data[430] ^ data[432] ^ data[433] ^ data[434] ^ data[435] ^ data[440] ^ data[441] ^ data[442] ^ data[443] ^ data[445] ^ data[447] ^ data[448] ^ data[450] ^ data[452] ^ data[455] ^ data[458] ^ data[459] ^ data[460] ^ data[462] ^ data[465] ^ data[467] ^ data[468] ^ data[469] ^ data[470] ^ data[472] ^ data[473] ^ data[474] ^ data[495];

assign temp_checkbits1[15] =   data[257] ^ data[258] ^ data[259] ^ data[260] ^ data[262] ^ data[263] ^ data[264] ^ data[267] ^ data[270] ^ data[271] ^ data[272] ^ data[275] ^ data[278] ^ data[280] ^ data[283] ^ data[284] ^ data[285] ^ data[287] ^ data[290] ^ data[292] ^ data[293] ^ data[296] ^ data[297] ^ data[301] ^ data[302] ^ data[304] ^ data[305] ^ data[309] ^ data[310] ^ data[312] ^ data[314] ^ data[315] ^ data[316] ^ data[317] ^ data[319] ^ data[320] ^ data[323] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[331] ^ data[332] ^ data[334] ^ data[335] ^ data[339] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[351] ^ data[352] ^ data[355] ^ data[356] ^ data[357] ^ data[360] ^ data[364] ^ data[365] ^ data[366] ^ data[367] ^ data[368] ^ data[370] ^ data[373] ^ data[374] ^ data[378] ^ data[379] ^ data[382] ^ data[383] ^ data[384] ^ data[385] ^ data[387] ^ data[392] ^ data[394] ^ data[398] ^ data[402] ^ data[403] ^ data[404] ^ data[405] ^ data[407] ^ data[409] ^ data[410] ^ data[412] ^ data[414] ^ data[415] ^ data[420] ^ data[421] ^ data[422] ^ data[423] ^ data[426] ^ data[427] ^ data[431] ^ data[433] ^ data[434] ^ data[435] ^ data[436] ^ data[441] ^ data[442] ^ data[443] ^ data[444] ^ data[446] ^ data[448] ^ data[449] ^ data[451] ^ data[453] ^ data[456] ^ data[459] ^ data[460] ^ data[461] ^ data[463] ^ data[466] ^ data[468] ^ data[469] ^ data[470] ^ data[471] ^ data[473] ^ data[474] ^ data[475] ^ data[496];

assign temp_checkbits1[14] =   data[257] ^ data[260] ^ data[261] ^ data[262] ^ data[264] ^ data[267] ^ data[271] ^ data[274] ^ data[277] ^ data[278] ^ data[279] ^ data[281] ^ data[282] ^ data[284] ^ data[286] ^ data[287] ^ data[297] ^ data[299] ^ data[300] ^ data[304] ^ data[308] ^ data[312] ^ data[313] ^ data[316] ^ data[317] ^ data[318] ^ data[323] ^ data[325] ^ data[328] ^ data[331] ^ data[332] ^ data[333] ^ data[336] ^ data[338] ^ data[340] ^ data[342] ^ data[345] ^ data[347] ^ data[348] ^ data[349] ^ data[351] ^ data[352] ^ data[353] ^ data[355] ^ data[361] ^ data[364] ^ data[365] ^ data[366] ^ data[367] ^ data[368] ^ data[371] ^ data[372] ^ data[373] ^ data[375] ^ data[376] ^ data[378] ^ data[381] ^ data[382] ^ data[384] ^ data[387] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[394] ^ data[396] ^ data[398] ^ data[403] ^ data[404] ^ data[406] ^ data[408] ^ data[412] ^ data[413] ^ data[414] ^ data[415] ^ data[416] ^ data[418] ^ data[420] ^ data[421] ^ data[422] ^ data[426] ^ data[427] ^ data[428] ^ data[432] ^ data[433] ^ data[434] ^ data[437] ^ data[443] ^ data[445] ^ data[446] ^ data[449] ^ data[453] ^ data[455] ^ data[457] ^ data[464] ^ data[466] ^ data[467] ^ data[468] ^ data[469] ^ data[470] ^ data[475] ^ data[497];

assign temp_checkbits1[13] =   data[256] ^ data[257] ^ data[259] ^ data[261] ^ data[267] ^ data[273] ^ data[274] ^ data[275] ^ data[276] ^ data[277] ^ data[279] ^ data[280] ^ data[283] ^ data[291] ^ data[293] ^ data[294] ^ data[299] ^ data[301] ^ data[302] ^ data[303] ^ data[304] ^ data[306] ^ data[308] ^ data[309] ^ data[310] ^ data[311] ^ data[312] ^ data[313] ^ data[314] ^ data[315] ^ data[317] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[323] ^ data[327] ^ data[330] ^ data[332] ^ data[333] ^ data[334] ^ data[335] ^ data[337] ^ data[338] ^ data[339] ^ data[341] ^ data[342] ^ data[343] ^ data[348] ^ data[350] ^ data[351] ^ data[352] ^ data[353] ^ data[354] ^ data[355] ^ data[357] ^ data[358] ^ data[362] ^ data[364] ^ data[365] ^ data[366] ^ data[367] ^ data[368] ^ data[377] ^ data[378] ^ data[380] ^ data[381] ^ data[386] ^ data[387] ^ data[388] ^ data[394] ^ data[396] ^ data[397] ^ data[398] ^ data[404] ^ data[407] ^ data[409] ^ data[410] ^ data[411] ^ data[412] ^ data[413] ^ data[415] ^ data[416] ^ data[417] ^ data[418] ^ data[419] ^ data[420] ^ data[421] ^ data[422] ^ data[424] ^ data[426] ^ data[427] ^ data[428] ^ data[429] ^ data[434] ^ data[436] ^ data[438] ^ data[442] ^ data[452] ^ data[453] ^ data[455] ^ data[456] ^ data[458] ^ data[460] ^ data[461] ^ data[462] ^ data[465] ^ data[466] ^ data[467] ^ data[469] ^ data[470] ^ data[472] ^ data[474] ^ data[498];

assign temp_checkbits1[12] =   data[256] ^ data[257] ^ data[258] ^ data[260] ^ data[262] ^ data[268] ^ data[274] ^ data[275] ^ data[276] ^ data[277] ^ data[278] ^ data[280] ^ data[281] ^ data[284] ^ data[292] ^ data[294] ^ data[295] ^ data[300] ^ data[302] ^ data[303] ^ data[304] ^ data[305] ^ data[307] ^ data[309] ^ data[310] ^ data[311] ^ data[312] ^ data[313] ^ data[314] ^ data[315] ^ data[316] ^ data[318] ^ data[319] ^ data[320] ^ data[321] ^ data[322] ^ data[324] ^ data[328] ^ data[331] ^ data[333] ^ data[334] ^ data[335] ^ data[336] ^ data[338] ^ data[339] ^ data[340] ^ data[342] ^ data[343] ^ data[344] ^ data[349] ^ data[351] ^ data[352] ^ data[353] ^ data[354] ^ data[355] ^ data[356] ^ data[358] ^ data[359] ^ data[363] ^ data[365] ^ data[366] ^ data[367] ^ data[368] ^ data[369] ^ data[378] ^ data[379] ^ data[381] ^ data[382] ^ data[387] ^ data[388] ^ data[389] ^ data[395] ^ data[397] ^ data[398] ^ data[399] ^ data[405] ^ data[408] ^ data[410] ^ data[411] ^ data[412] ^ data[413] ^ data[414] ^ data[416] ^ data[417] ^ data[418] ^ data[419] ^ data[420] ^ data[421] ^ data[422] ^ data[423] ^ data[425] ^ data[427] ^ data[428] ^ data[429] ^ data[430] ^ data[435] ^ data[437] ^ data[439] ^ data[443] ^ data[453] ^ data[454] ^ data[456] ^ data[457] ^ data[459] ^ data[461] ^ data[462] ^ data[463] ^ data[466] ^ data[467] ^ data[468] ^ data[470] ^ data[471] ^ data[473] ^ data[475] ^ data[499];

assign temp_checkbits1[11] =   data[256] ^ data[261] ^ data[262] ^ data[265] ^ data[267] ^ data[268] ^ data[269] ^ data[272] ^ data[273] ^ data[274] ^ data[275] ^ data[279] ^ data[281] ^ data[287] ^ data[288] ^ data[291] ^ data[294] ^ data[295] ^ data[296] ^ data[298] ^ data[299] ^ data[300] ^ data[301] ^ data[302] ^ data[313] ^ data[314] ^ data[316] ^ data[317] ^ data[319] ^ data[322] ^ data[324] ^ data[325] ^ data[326] ^ data[327] ^ data[330] ^ data[332] ^ data[334] ^ data[336] ^ data[337] ^ data[338] ^ data[339] ^ data[340] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[349] ^ data[350] ^ data[351] ^ data[352] ^ data[353] ^ data[354] ^ data[358] ^ data[359] ^ data[360] ^ data[366] ^ data[367] ^ data[368] ^ data[370] ^ data[372] ^ data[373] ^ data[374] ^ data[376] ^ data[378] ^ data[381] ^ data[385] ^ data[386] ^ data[387] ^ data[388] ^ data[391] ^ data[392] ^ data[393] ^ data[394] ^ data[395] ^ data[400] ^ data[405] ^ data[406] ^ data[409] ^ data[410] ^ data[413] ^ data[415] ^ data[417] ^ data[419] ^ data[421] ^ data[422] ^ data[428] ^ data[429] ^ data[430] ^ data[431] ^ data[433] ^ data[435] ^ data[438] ^ data[440] ^ data[442] ^ data[446] ^ data[447] ^ data[450] ^ data[452] ^ data[453] ^ data[457] ^ data[458] ^ data[461] ^ data[463] ^ data[464] ^ data[466] ^ data[467] ^ data[469] ^ data[500];

assign temp_checkbits1[10] =   data[256] ^ data[257] ^ data[262] ^ data[263] ^ data[266] ^ data[268] ^ data[269] ^ data[270] ^ data[273] ^ data[274] ^ data[275] ^ data[276] ^ data[280] ^ data[282] ^ data[288] ^ data[289] ^ data[292] ^ data[295] ^ data[296] ^ data[297] ^ data[299] ^ data[300] ^ data[301] ^ data[302] ^ data[303] ^ data[314] ^ data[315] ^ data[317] ^ data[318] ^ data[320] ^ data[323] ^ data[325] ^ data[326] ^ data[327] ^ data[328] ^ data[331] ^ data[333] ^ data[335] ^ data[337] ^ data[338] ^ data[339] ^ data[340] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[350] ^ data[351] ^ data[352] ^ data[353] ^ data[354] ^ data[355] ^ data[359] ^ data[360] ^ data[361] ^ data[367] ^ data[368] ^ data[369] ^ data[371] ^ data[373] ^ data[374] ^ data[375] ^ data[377] ^ data[379] ^ data[382] ^ data[386] ^ data[387] ^ data[388] ^ data[389] ^ data[392] ^ data[393] ^ data[394] ^ data[395] ^ data[396] ^ data[401] ^ data[406] ^ data[407] ^ data[410] ^ data[411] ^ data[414] ^ data[416] ^ data[418] ^ data[420] ^ data[422] ^ data[423] ^ data[429] ^ data[430] ^ data[431] ^ data[432] ^ data[434] ^ data[436] ^ data[439] ^ data[441] ^ data[443] ^ data[447] ^ data[448] ^ data[451] ^ data[453] ^ data[454] ^ data[458] ^ data[459] ^ data[462] ^ data[464] ^ data[465] ^ data[467] ^ data[468] ^ data[470] ^ data[501];

assign temp_checkbits1[9] =   data[256] ^ data[257] ^ data[258] ^ data[263] ^ data[264] ^ data[267] ^ data[269] ^ data[270] ^ data[271] ^ data[274] ^ data[275] ^ data[276] ^ data[277] ^ data[281] ^ data[283] ^ data[289] ^ data[290] ^ data[293] ^ data[296] ^ data[297] ^ data[298] ^ data[300] ^ data[301] ^ data[302] ^ data[303] ^ data[304] ^ data[315] ^ data[316] ^ data[318] ^ data[319] ^ data[321] ^ data[324] ^ data[326] ^ data[327] ^ data[328] ^ data[329] ^ data[332] ^ data[334] ^ data[336] ^ data[338] ^ data[339] ^ data[340] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[348] ^ data[351] ^ data[352] ^ data[353] ^ data[354] ^ data[355] ^ data[356] ^ data[360] ^ data[361] ^ data[362] ^ data[368] ^ data[369] ^ data[370] ^ data[372] ^ data[374] ^ data[375] ^ data[376] ^ data[378] ^ data[380] ^ data[383] ^ data[387] ^ data[388] ^ data[389] ^ data[390] ^ data[393] ^ data[394] ^ data[395] ^ data[396] ^ data[397] ^ data[402] ^ data[407] ^ data[408] ^ data[411] ^ data[412] ^ data[415] ^ data[417] ^ data[419] ^ data[421] ^ data[423] ^ data[424] ^ data[430] ^ data[431] ^ data[432] ^ data[433] ^ data[435] ^ data[437] ^ data[440] ^ data[442] ^ data[444] ^ data[448] ^ data[449] ^ data[452] ^ data[454] ^ data[455] ^ data[459] ^ data[460] ^ data[463] ^ data[465] ^ data[466] ^ data[468] ^ data[469] ^ data[471] ^ data[502];

assign temp_checkbits1[8] =   data[257] ^ data[258] ^ data[259] ^ data[264] ^ data[265] ^ data[268] ^ data[270] ^ data[271] ^ data[272] ^ data[275] ^ data[276] ^ data[277] ^ data[278] ^ data[282] ^ data[284] ^ data[290] ^ data[291] ^ data[294] ^ data[297] ^ data[298] ^ data[299] ^ data[301] ^ data[302] ^ data[303] ^ data[304] ^ data[305] ^ data[316] ^ data[317] ^ data[319] ^ data[320] ^ data[322] ^ data[325] ^ data[327] ^ data[328] ^ data[329] ^ data[330] ^ data[333] ^ data[335] ^ data[337] ^ data[339] ^ data[340] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[348] ^ data[349] ^ data[352] ^ data[353] ^ data[354] ^ data[355] ^ data[356] ^ data[357] ^ data[361] ^ data[362] ^ data[363] ^ data[369] ^ data[370] ^ data[371] ^ data[373] ^ data[375] ^ data[376] ^ data[377] ^ data[379] ^ data[381] ^ data[384] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[394] ^ data[395] ^ data[396] ^ data[397] ^ data[398] ^ data[403] ^ data[408] ^ data[409] ^ data[412] ^ data[413] ^ data[416] ^ data[418] ^ data[420] ^ data[422] ^ data[424] ^ data[425] ^ data[431] ^ data[432] ^ data[433] ^ data[434] ^ data[436] ^ data[438] ^ data[441] ^ data[443] ^ data[445] ^ data[449] ^ data[450] ^ data[453] ^ data[455] ^ data[456] ^ data[460] ^ data[461] ^ data[464] ^ data[466] ^ data[467] ^ data[469] ^ data[470] ^ data[472] ^ data[503];

assign temp_checkbits1[7] =   data[256] ^ data[258] ^ data[259] ^ data[260] ^ data[265] ^ data[266] ^ data[269] ^ data[271] ^ data[272] ^ data[273] ^ data[276] ^ data[277] ^ data[278] ^ data[279] ^ data[283] ^ data[285] ^ data[291] ^ data[292] ^ data[295] ^ data[298] ^ data[299] ^ data[300] ^ data[302] ^ data[303] ^ data[304] ^ data[305] ^ data[306] ^ data[317] ^ data[318] ^ data[320] ^ data[321] ^ data[323] ^ data[326] ^ data[328] ^ data[329] ^ data[330] ^ data[331] ^ data[334] ^ data[336] ^ data[338] ^ data[340] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[348] ^ data[349] ^ data[350] ^ data[353] ^ data[354] ^ data[355] ^ data[356] ^ data[357] ^ data[358] ^ data[362] ^ data[363] ^ data[364] ^ data[370] ^ data[371] ^ data[372] ^ data[374] ^ data[376] ^ data[377] ^ data[378] ^ data[380] ^ data[382] ^ data[385] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[395] ^ data[396] ^ data[397] ^ data[398] ^ data[399] ^ data[404] ^ data[409] ^ data[410] ^ data[413] ^ data[414] ^ data[417] ^ data[419] ^ data[421] ^ data[423] ^ data[425] ^ data[426] ^ data[432] ^ data[433] ^ data[434] ^ data[435] ^ data[437] ^ data[439] ^ data[442] ^ data[444] ^ data[446] ^ data[450] ^ data[451] ^ data[454] ^ data[456] ^ data[457] ^ data[461] ^ data[462] ^ data[465] ^ data[467] ^ data[468] ^ data[470] ^ data[471] ^ data[473] ^ data[504];

assign temp_checkbits1[6] =   data[256] ^ data[257] ^ data[259] ^ data[260] ^ data[261] ^ data[266] ^ data[267] ^ data[270] ^ data[272] ^ data[273] ^ data[274] ^ data[277] ^ data[278] ^ data[279] ^ data[280] ^ data[284] ^ data[286] ^ data[292] ^ data[293] ^ data[296] ^ data[299] ^ data[300] ^ data[301] ^ data[303] ^ data[304] ^ data[305] ^ data[306] ^ data[307] ^ data[318] ^ data[319] ^ data[321] ^ data[322] ^ data[324] ^ data[327] ^ data[329] ^ data[330] ^ data[331] ^ data[332] ^ data[335] ^ data[337] ^ data[339] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[348] ^ data[349] ^ data[350] ^ data[351] ^ data[354] ^ data[355] ^ data[356] ^ data[357] ^ data[358] ^ data[359] ^ data[363] ^ data[364] ^ data[365] ^ data[371] ^ data[372] ^ data[373] ^ data[375] ^ data[377] ^ data[378] ^ data[379] ^ data[381] ^ data[383] ^ data[386] ^ data[390] ^ data[391] ^ data[392] ^ data[393] ^ data[396] ^ data[397] ^ data[398] ^ data[399] ^ data[400] ^ data[405] ^ data[410] ^ data[411] ^ data[414] ^ data[415] ^ data[418] ^ data[420] ^ data[422] ^ data[424] ^ data[426] ^ data[427] ^ data[433] ^ data[434] ^ data[435] ^ data[436] ^ data[438] ^ data[440] ^ data[443] ^ data[445] ^ data[447] ^ data[451] ^ data[452] ^ data[455] ^ data[457] ^ data[458] ^ data[462] ^ data[463] ^ data[466] ^ data[468] ^ data[469] ^ data[471] ^ data[472] ^ data[474] ^ data[505];

assign temp_checkbits1[5] =   data[257] ^ data[258] ^ data[260] ^ data[261] ^ data[262] ^ data[267] ^ data[268] ^ data[271] ^ data[273] ^ data[274] ^ data[275] ^ data[278] ^ data[279] ^ data[280] ^ data[281] ^ data[285] ^ data[287] ^ data[293] ^ data[294] ^ data[297] ^ data[300] ^ data[301] ^ data[302] ^ data[304] ^ data[305] ^ data[306] ^ data[307] ^ data[308] ^ data[319] ^ data[320] ^ data[322] ^ data[323] ^ data[325] ^ data[328] ^ data[330] ^ data[331] ^ data[332] ^ data[333] ^ data[336] ^ data[338] ^ data[340] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[348] ^ data[349] ^ data[350] ^ data[351] ^ data[352] ^ data[355] ^ data[356] ^ data[357] ^ data[358] ^ data[359] ^ data[360] ^ data[364] ^ data[365] ^ data[366] ^ data[372] ^ data[373] ^ data[374] ^ data[376] ^ data[378] ^ data[379] ^ data[380] ^ data[382] ^ data[384] ^ data[387] ^ data[391] ^ data[392] ^ data[393] ^ data[394] ^ data[397] ^ data[398] ^ data[399] ^ data[400] ^ data[401] ^ data[406] ^ data[411] ^ data[412] ^ data[415] ^ data[416] ^ data[419] ^ data[421] ^ data[423] ^ data[425] ^ data[427] ^ data[428] ^ data[434] ^ data[435] ^ data[436] ^ data[437] ^ data[439] ^ data[441] ^ data[444] ^ data[446] ^ data[448] ^ data[452] ^ data[453] ^ data[456] ^ data[458] ^ data[459] ^ data[463] ^ data[464] ^ data[467] ^ data[469] ^ data[470] ^ data[472] ^ data[473] ^ data[475] ^ data[506];

assign temp_checkbits1[4] =   data[256] ^ data[257] ^ data[261] ^ data[265] ^ data[267] ^ data[269] ^ data[273] ^ data[275] ^ data[277] ^ data[278] ^ data[279] ^ data[280] ^ data[281] ^ data[285] ^ data[286] ^ data[287] ^ data[291] ^ data[293] ^ data[295] ^ data[299] ^ data[300] ^ data[301] ^ data[304] ^ data[307] ^ data[309] ^ data[310] ^ data[311] ^ data[312] ^ data[315] ^ data[327] ^ data[330] ^ data[331] ^ data[332] ^ data[333] ^ data[334] ^ data[335] ^ data[337] ^ data[338] ^ data[339] ^ data[341] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[347] ^ data[348] ^ data[350] ^ data[352] ^ data[353] ^ data[355] ^ data[359] ^ data[360] ^ data[361] ^ data[364] ^ data[365] ^ data[366] ^ data[367] ^ data[369] ^ data[372] ^ data[375] ^ data[376] ^ data[377] ^ data[378] ^ data[382] ^ data[386] ^ data[387] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[396] ^ data[400] ^ data[401] ^ data[402] ^ data[405] ^ data[407] ^ data[410] ^ data[411] ^ data[413] ^ data[414] ^ data[416] ^ data[417] ^ data[418] ^ data[422] ^ data[423] ^ data[428] ^ data[429] ^ data[433] ^ data[437] ^ data[438] ^ data[440] ^ data[444] ^ data[445] ^ data[446] ^ data[449] ^ data[450] ^ data[452] ^ data[455] ^ data[457] ^ data[459] ^ data[461] ^ data[462] ^ data[464] ^ data[465] ^ data[466] ^ data[470] ^ data[472] ^ data[473] ^ data[507];

assign temp_checkbits1[3] =   data[257] ^ data[258] ^ data[262] ^ data[266] ^ data[268] ^ data[270] ^ data[274] ^ data[276] ^ data[278] ^ data[279] ^ data[280] ^ data[281] ^ data[282] ^ data[286] ^ data[287] ^ data[288] ^ data[292] ^ data[294] ^ data[296] ^ data[300] ^ data[301] ^ data[302] ^ data[305] ^ data[308] ^ data[310] ^ data[311] ^ data[312] ^ data[313] ^ data[316] ^ data[328] ^ data[331] ^ data[332] ^ data[333] ^ data[334] ^ data[335] ^ data[336] ^ data[338] ^ data[339] ^ data[340] ^ data[342] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[348] ^ data[349] ^ data[351] ^ data[353] ^ data[354] ^ data[356] ^ data[360] ^ data[361] ^ data[362] ^ data[365] ^ data[366] ^ data[367] ^ data[368] ^ data[370] ^ data[373] ^ data[376] ^ data[377] ^ data[378] ^ data[379] ^ data[383] ^ data[387] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[397] ^ data[401] ^ data[402] ^ data[403] ^ data[406] ^ data[408] ^ data[411] ^ data[412] ^ data[414] ^ data[415] ^ data[417] ^ data[418] ^ data[419] ^ data[423] ^ data[424] ^ data[429] ^ data[430] ^ data[434] ^ data[438] ^ data[439] ^ data[441] ^ data[445] ^ data[446] ^ data[447] ^ data[450] ^ data[451] ^ data[453] ^ data[456] ^ data[458] ^ data[460] ^ data[462] ^ data[463] ^ data[465] ^ data[466] ^ data[467] ^ data[471] ^ data[473] ^ data[474] ^ data[508];

assign temp_checkbits1[2] =   data[256] ^ data[258] ^ data[259] ^ data[263] ^ data[267] ^ data[269] ^ data[271] ^ data[275] ^ data[277] ^ data[279] ^ data[280] ^ data[281] ^ data[282] ^ data[283] ^ data[287] ^ data[288] ^ data[289] ^ data[293] ^ data[295] ^ data[297] ^ data[301] ^ data[302] ^ data[303] ^ data[306] ^ data[309] ^ data[311] ^ data[312] ^ data[313] ^ data[314] ^ data[317] ^ data[329] ^ data[332] ^ data[333] ^ data[334] ^ data[335] ^ data[336] ^ data[337] ^ data[339] ^ data[340] ^ data[341] ^ data[343] ^ data[344] ^ data[345] ^ data[346] ^ data[347] ^ data[349] ^ data[350] ^ data[352] ^ data[354] ^ data[355] ^ data[357] ^ data[361] ^ data[362] ^ data[363] ^ data[366] ^ data[367] ^ data[368] ^ data[369] ^ data[371] ^ data[374] ^ data[377] ^ data[378] ^ data[379] ^ data[380] ^ data[384] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[393] ^ data[398] ^ data[402] ^ data[403] ^ data[404] ^ data[407] ^ data[409] ^ data[412] ^ data[413] ^ data[415] ^ data[416] ^ data[418] ^ data[419] ^ data[420] ^ data[424] ^ data[425] ^ data[430] ^ data[431] ^ data[435] ^ data[439] ^ data[440] ^ data[442] ^ data[446] ^ data[447] ^ data[448] ^ data[451] ^ data[452] ^ data[454] ^ data[457] ^ data[459] ^ data[461] ^ data[463] ^ data[464] ^ data[466] ^ data[467] ^ data[468] ^ data[472] ^ data[474] ^ data[475] ^ data[509];

assign temp_checkbits1[1] =   data[258] ^ data[260] ^ data[262] ^ data[263] ^ data[264] ^ data[265] ^ data[267] ^ data[270] ^ data[273] ^ data[274] ^ data[277] ^ data[280] ^ data[281] ^ data[283] ^ data[284] ^ data[285] ^ data[287] ^ data[289] ^ data[290] ^ data[291] ^ data[293] ^ data[296] ^ data[299] ^ data[300] ^ data[305] ^ data[306] ^ data[307] ^ data[308] ^ data[311] ^ data[313] ^ data[314] ^ data[318] ^ data[320] ^ data[321] ^ data[323] ^ data[324] ^ data[326] ^ data[327] ^ data[329] ^ data[333] ^ data[334] ^ data[336] ^ data[337] ^ data[340] ^ data[341] ^ data[344] ^ data[345] ^ data[347] ^ data[348] ^ data[349] ^ data[350] ^ data[353] ^ data[357] ^ data[362] ^ data[363] ^ data[367] ^ data[368] ^ data[370] ^ data[373] ^ data[374] ^ data[375] ^ data[376] ^ data[382] ^ data[383] ^ data[386] ^ data[387] ^ data[395] ^ data[396] ^ data[398] ^ data[403] ^ data[404] ^ data[408] ^ data[411] ^ data[412] ^ data[413] ^ data[416] ^ data[417] ^ data[418] ^ data[419] ^ data[421] ^ data[423] ^ data[424] ^ data[425] ^ data[431] ^ data[432] ^ data[433] ^ data[435] ^ data[440] ^ data[441] ^ data[442] ^ data[443] ^ data[444] ^ data[446] ^ data[448] ^ data[449] ^ data[450] ^ data[454] ^ data[458] ^ data[461] ^ data[464] ^ data[465] ^ data[466] ^ data[467] ^ data[469] ^ data[471] ^ data[472] ^ data[473] ^ data[474] ^ data[475] ^ data[510];

assign temp_checkbits1[0] =   data[256] ^ data[257] ^ data[258] ^ data[261] ^ data[262] ^ data[264] ^ data[266] ^ data[267] ^ data[271] ^ data[272] ^ data[273] ^ data[275] ^ data[276] ^ data[277] ^ data[281] ^ data[284] ^ data[286] ^ data[287] ^ data[290] ^ data[292] ^ data[293] ^ data[297] ^ data[298] ^ data[299] ^ data[301] ^ data[302] ^ data[303] ^ data[304] ^ data[305] ^ data[307] ^ data[309] ^ data[310] ^ data[311] ^ data[314] ^ data[319] ^ data[320] ^ data[322] ^ data[323] ^ data[325] ^ data[326] ^ data[328] ^ data[329] ^ data[334] ^ data[337] ^ data[341] ^ data[345] ^ data[348] ^ data[350] ^ data[354] ^ data[355] ^ data[356] ^ data[357] ^ data[363] ^ data[368] ^ data[371] ^ data[372] ^ data[373] ^ data[375] ^ data[377] ^ data[378] ^ data[379] ^ data[380] ^ data[381] ^ data[382] ^ data[384] ^ data[385] ^ data[386] ^ data[388] ^ data[389] ^ data[390] ^ data[391] ^ data[392] ^ data[393] ^ data[394] ^ data[395] ^ data[397] ^ data[398] ^ data[404] ^ data[409] ^ data[410] ^ data[411] ^ data[413] ^ data[417] ^ data[419] ^ data[422] ^ data[423] ^ data[425] ^ data[432] ^ data[434] ^ data[435] ^ data[441] ^ data[443] ^ data[445] ^ data[446] ^ data[449] ^ data[451] ^ data[452] ^ data[453] ^ data[454] ^ data[459] ^ data[460] ^ data[461] ^ data[465] ^ data[467] ^ data[470] ^ data[471] ^ data[473] ^ data[475] ^ data[511];





   
assign    checkbits0_out = temp_checkbits0;
assign    checkbits1_out = temp_checkbits1;





   

endmodule //-- ocx_dlx_crc
